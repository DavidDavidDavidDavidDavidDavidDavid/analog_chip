magic
tech sky130A
magscale 1 2
timestamp 1685060018
<< nwell >>
rect 5326 749 6141 1070
rect 6698 824 6760 978
rect 5322 -491 5875 -170
rect 6642 -224 6846 -90
rect 6710 -278 6722 -272
rect 6772 -278 6774 -276
rect 6710 -386 6720 -278
rect 6710 -398 6774 -386
rect 5320 -1291 5872 -970
rect 6624 -1018 6856 -906
rect 6662 -1020 6816 -1018
rect 6648 -1820 6856 -1714
rect 6652 -2604 6874 -2500
rect 6652 -3396 6874 -3292
rect 6640 -4222 6862 -4118
rect 6618 -5028 6840 -4924
rect 6622 -5844 6856 -5710
rect 6638 -7006 6860 -6902
<< pwell >>
rect 5701 483 7740 691
rect 6640 424 6848 483
rect 5296 -757 8183 -549
rect 6654 -822 6862 -757
rect 5292 -1557 8222 -1349
rect 6644 -1614 6852 -1557
rect 5331 -2357 8168 -2149
rect 6648 -2422 6856 -2357
rect 5299 -3159 8204 -2949
rect 6640 -3226 6848 -3159
rect 5324 -3963 8183 -3749
rect 6636 -4032 6844 -3963
rect 5323 -4757 8203 -4549
rect 6654 -4818 6862 -4757
rect 5296 -5557 8195 -5349
rect 6648 -5608 6856 -5557
rect 5326 -6367 8196 -6149
rect 6632 -6428 6840 -6367
rect 6507 -7334 6965 -7330
rect 5739 -7542 7732 -7334
rect 6646 -7594 6854 -7542
<< psubdiff >>
rect 6676 440 6700 474
rect 6750 440 6774 474
rect 6698 -800 6722 -766
rect 6772 -800 6796 -766
rect 6696 -1600 6720 -1566
rect 6770 -1600 6794 -1566
rect 6698 -2400 6722 -2366
rect 6772 -2400 6796 -2366
rect 6698 -3200 6722 -3166
rect 6772 -3200 6796 -3166
rect 6698 -4000 6722 -3966
rect 6772 -4000 6796 -3966
rect 6698 -4800 6722 -4766
rect 6772 -4800 6796 -4766
rect 6698 -5600 6722 -5566
rect 6772 -5600 6796 -5566
rect 6698 -6400 6722 -6366
rect 6772 -6400 6796 -6366
rect 6698 -7582 6722 -7548
rect 6772 -7582 6796 -7548
<< nsubdiff >>
rect 6704 938 6750 962
rect 6704 842 6750 866
rect 6696 -194 6720 -160
rect 6770 -194 6794 -160
rect 6700 -994 6724 -960
rect 6774 -994 6798 -960
rect 6700 -1794 6724 -1760
rect 6774 -1794 6798 -1760
rect 6698 -2592 6722 -2558
rect 6772 -2592 6796 -2558
rect 6698 -3394 6722 -3360
rect 6772 -3394 6796 -3360
rect 6700 -4194 6724 -4160
rect 6774 -4194 6798 -4160
rect 6700 -4994 6724 -4960
rect 6774 -4994 6798 -4960
rect 6698 -5794 6722 -5760
rect 6772 -5794 6796 -5760
rect 6700 -6982 6724 -6948
rect 6774 -6982 6798 -6948
<< psubdiffcont >>
rect 6700 440 6750 474
rect 6722 -800 6772 -766
rect 6720 -1600 6770 -1566
rect 6722 -2400 6772 -2366
rect 6722 -3200 6772 -3166
rect 6722 -4000 6772 -3966
rect 6722 -4800 6772 -4766
rect 6722 -5600 6772 -5566
rect 6722 -6400 6772 -6366
rect 6722 -7582 6772 -7548
<< nsubdiffcont >>
rect 6704 866 6750 938
rect 6720 -194 6770 -160
rect 6724 -994 6774 -960
rect 6724 -1794 6774 -1760
rect 6722 -2592 6772 -2558
rect 6722 -3394 6772 -3360
rect 6724 -4194 6774 -4160
rect 6724 -4994 6774 -4960
rect 6722 -5794 6772 -5760
rect 6724 -6982 6774 -6948
<< locali >>
rect 5713 935 5757 1047
rect 6565 1015 6815 1049
rect 6704 938 6750 1015
rect 7693 935 7737 1038
rect 6704 850 6750 866
rect 5707 483 5765 599
rect 6565 474 6855 505
rect 7683 486 7741 599
rect 6565 471 6700 474
rect 6684 440 6700 471
rect 6750 471 6855 474
rect 6750 440 6766 471
rect 6704 -191 6720 -160
rect 6589 -194 6720 -191
rect 6770 -191 6786 -160
rect 6770 -194 6903 -191
rect 5294 -305 5338 -195
rect 6589 -225 6903 -194
rect 8157 -305 8201 -202
rect 5559 -493 5609 -489
rect 5559 -571 5609 -543
rect 7903 -587 7953 -543
rect 5287 -750 5345 -641
rect 6593 -766 6957 -735
rect 8151 -757 8209 -641
rect 6593 -769 6722 -766
rect 6706 -800 6722 -769
rect 6772 -769 6957 -766
rect 6772 -800 6788 -769
rect 6708 -991 6724 -960
rect 6589 -994 6724 -991
rect 6774 -991 6790 -960
rect 6774 -994 6947 -991
rect 5299 -1105 5343 -994
rect 6589 -1025 6947 -994
rect 8158 -1105 8202 -1000
rect 5560 -1282 5610 -1278
rect 5560 -1360 5610 -1332
rect 7903 -1373 7953 -1327
rect 5287 -1554 5345 -1441
rect 6595 -1566 6883 -1535
rect 8151 -1564 8209 -1441
rect 6595 -1569 6720 -1566
rect 6704 -1600 6720 -1569
rect 6770 -1569 6883 -1566
rect 6770 -1600 6786 -1569
rect 6708 -1791 6724 -1760
rect 6589 -1794 6724 -1791
rect 6774 -1791 6790 -1760
rect 6774 -1794 6881 -1791
rect 5298 -1905 5342 -1804
rect 6589 -1825 6881 -1794
rect 8156 -1905 8200 -1795
rect 5560 -2082 5610 -2078
rect 5560 -2160 5610 -2132
rect 7903 -2169 7953 -2125
rect 5287 -2365 5345 -2241
rect 6601 -2366 6911 -2335
rect 8151 -2359 8209 -2241
rect 6601 -2369 6722 -2366
rect 6706 -2400 6722 -2369
rect 6772 -2369 6911 -2366
rect 6772 -2400 6788 -2369
rect 6706 -2591 6722 -2558
rect 5293 -2789 5343 -2591
rect 6589 -2592 6722 -2591
rect 6772 -2591 6788 -2558
rect 6772 -2592 6907 -2591
rect 6589 -2625 6907 -2592
rect 8160 -2705 8204 -2602
rect 5560 -2882 5610 -2878
rect 5560 -2960 5610 -2932
rect 7903 -2971 7953 -2933
rect 5287 -3169 5345 -3041
rect 6609 -3166 6879 -3135
rect 8151 -3163 8209 -3041
rect 6609 -3169 6722 -3166
rect 6706 -3200 6722 -3169
rect 6772 -3169 6879 -3166
rect 6772 -3200 6788 -3169
rect 6706 -3391 6722 -3360
rect 6589 -3394 6722 -3391
rect 6772 -3391 6788 -3360
rect 6772 -3394 6923 -3391
rect 5294 -3505 5338 -3399
rect 6589 -3425 6923 -3394
rect 8159 -3505 8203 -3398
rect 5560 -3678 5610 -3674
rect 5560 -3756 5610 -3728
rect 7903 -3773 7953 -3731
rect 5287 -3954 5345 -3841
rect 6595 -3966 6875 -3935
rect 8151 -3966 8209 -3841
rect 6595 -3969 6722 -3966
rect 6706 -4000 6722 -3969
rect 6772 -3969 6875 -3966
rect 6772 -4000 6788 -3969
rect 6708 -4191 6724 -4160
rect 6589 -4194 6724 -4191
rect 6774 -4191 6790 -4160
rect 6774 -4194 6895 -4191
rect 5298 -4305 5342 -4196
rect 6589 -4225 6895 -4194
rect 8158 -4305 8202 -4203
rect 5560 -4474 5610 -4470
rect 5560 -4552 5610 -4524
rect 7903 -4561 7953 -4527
rect 5287 -4762 5345 -4641
rect 6589 -4766 6889 -4735
rect 8151 -4766 8209 -4641
rect 6589 -4769 6722 -4766
rect 6706 -4800 6722 -4769
rect 6772 -4769 6889 -4766
rect 6772 -4800 6788 -4769
rect 6708 -4991 6724 -4960
rect 6589 -4994 6724 -4991
rect 6774 -4991 6790 -4960
rect 6774 -4994 6913 -4991
rect 5294 -5105 5338 -5009
rect 6589 -5025 6913 -4994
rect 8154 -5105 8198 -4998
rect 5560 -5276 5610 -5272
rect 5560 -5354 5610 -5326
rect 7903 -5369 7953 -5327
rect 5287 -5559 5345 -5441
rect 6613 -5566 6877 -5535
rect 8151 -5558 8209 -5441
rect 6613 -5569 6722 -5566
rect 6706 -5600 6722 -5569
rect 6772 -5569 6877 -5566
rect 6772 -5600 6788 -5569
rect 6706 -5791 6722 -5760
rect 6589 -5794 6722 -5791
rect 6772 -5791 6788 -5760
rect 6772 -5794 6891 -5791
rect 5296 -5905 5340 -5799
rect 6589 -5825 6891 -5794
rect 8152 -5905 8196 -5796
rect 5560 -6070 5610 -6066
rect 5560 -6148 5610 -6120
rect 7903 -6165 7953 -6137
rect 5287 -6360 5345 -6241
rect 6535 -6366 6905 -6335
rect 8151 -6351 8209 -6241
rect 6535 -6369 6722 -6366
rect 6706 -6400 6722 -6369
rect 6772 -6369 6905 -6366
rect 6772 -6400 6788 -6369
rect 6708 -6972 6724 -6948
rect 6593 -6982 6724 -6972
rect 6774 -6972 6790 -6948
rect 6774 -6982 6875 -6972
rect 5738 -7086 5782 -6982
rect 6593 -7006 6875 -6982
rect 7716 -7086 7760 -6975
rect 5730 -7534 5788 -7422
rect 6611 -7548 6843 -7516
rect 7706 -7525 7764 -7422
rect 6611 -7550 6722 -7548
rect 6706 -7582 6722 -7550
rect 6772 -7550 6843 -7548
rect 6772 -7582 6788 -7550
<< viali >>
rect 5876 754 5946 814
rect 7504 760 7564 820
rect 6046 704 6086 744
rect 6176 704 6216 744
rect 6326 704 6366 744
rect 6456 704 6496 744
rect 6936 704 6976 744
rect 7066 704 7106 744
rect 7216 704 7256 744
rect 7346 704 7386 744
rect 5876 634 5946 694
rect 7503 631 7572 700
rect 5468 -533 5507 -494
rect 5559 -543 5609 -493
rect 7814 -533 7853 -494
rect 7903 -543 7953 -493
rect 5468 -1330 5507 -1291
rect 5560 -1332 5610 -1282
rect 7804 -1333 7843 -1294
rect 7903 -1327 7953 -1277
rect 5466 -2131 5505 -2092
rect 5560 -2132 5610 -2082
rect 7813 -2130 7852 -2091
rect 7903 -2125 7953 -2075
rect 5464 -2931 5503 -2892
rect 5560 -2932 5610 -2882
rect 7808 -2931 7847 -2892
rect 7903 -2933 7953 -2883
rect 5457 -3732 5496 -3693
rect 5560 -3728 5610 -3678
rect 7808 -3733 7847 -3694
rect 7903 -3731 7953 -3681
rect 5466 -4531 5505 -4492
rect 5560 -4524 5610 -4474
rect 7807 -4531 7846 -4492
rect 7903 -4527 7953 -4477
rect 5464 -5330 5503 -5291
rect 5560 -5326 5610 -5276
rect 7802 -5329 7841 -5290
rect 7903 -5327 7953 -5277
rect 5463 -6132 5502 -6093
rect 5560 -6120 5610 -6070
rect 7807 -6134 7846 -6095
rect 7903 -6137 7953 -6087
rect 6634 -7260 6694 -7200
rect 7534 -7260 7594 -7200
rect 6075 -7310 6115 -7270
rect 6205 -7310 6245 -7270
rect 6355 -7310 6395 -7270
rect 6485 -7310 6525 -7270
rect 6963 -7314 7003 -7274
rect 7093 -7314 7133 -7274
rect 7243 -7314 7283 -7274
rect 7373 -7314 7413 -7274
rect 6634 -7388 6694 -7328
rect 7534 -7388 7594 -7328
<< metal1 >>
rect 4768 1928 4828 1934
rect 5092 1930 5152 2270
rect 5320 2060 5380 2354
rect 5320 1990 5380 1996
rect 2776 1868 4768 1928
rect 4864 1870 4870 1930
rect 4930 1870 5152 1930
rect 2776 1750 2836 1868
rect 4768 1862 4828 1868
rect 7924 1866 7984 2264
rect 9218 1884 9278 2266
rect 7924 1806 7970 1866
rect 8030 1806 8036 1866
rect 8764 1824 8770 1884
rect 8830 1824 9278 1884
rect 8884 1602 8890 1662
rect 8950 1602 9390 1662
rect 5036 984 5042 1080
rect 5138 984 7786 1080
rect 5866 820 5876 824
rect 5864 754 5876 820
rect 5946 820 5956 824
rect 7492 820 7576 826
rect 5946 754 5958 820
rect 7492 760 7504 820
rect 7564 760 7576 820
rect 5864 748 5958 754
rect 6036 754 6096 760
rect 5864 694 5958 700
rect 6034 698 6036 750
rect 6166 754 6226 760
rect 3970 630 4650 690
rect 4710 630 4716 690
rect 5864 634 5876 694
rect 5946 634 5958 694
rect 6096 698 6098 750
rect 6164 698 6166 750
rect 6316 754 6376 760
rect 6036 688 6096 694
rect 6226 698 6228 750
rect 6314 698 6316 750
rect 6446 754 6506 760
rect 6166 688 6226 694
rect 6376 698 6378 750
rect 6444 698 6446 750
rect 6926 754 6986 760
rect 6316 688 6376 694
rect 6506 698 6508 750
rect 6924 698 6926 750
rect 7056 754 7116 760
rect 6446 688 6506 694
rect 6986 698 6988 750
rect 7054 698 7056 750
rect 7206 754 7266 760
rect 6926 688 6986 694
rect 7116 698 7118 750
rect 7204 698 7206 750
rect 7336 754 7396 760
rect 7492 754 7576 760
rect 7056 688 7116 694
rect 7266 698 7268 750
rect 7334 698 7336 750
rect 7206 688 7266 694
rect 7396 698 7398 750
rect 7491 700 7584 706
rect 7336 688 7396 694
rect 5864 628 5958 634
rect 7491 631 7503 700
rect 7572 631 7584 700
rect 7491 625 7584 631
rect 5500 440 8416 536
rect 8512 440 8518 536
rect 4530 310 4590 316
rect 2690 250 4530 310
rect 2690 50 2750 250
rect 4530 244 4590 250
rect 9010 196 9070 202
rect 11420 196 11480 550
rect 9070 136 11480 196
rect 9010 130 9070 136
rect 5056 -256 5062 -160
rect 5158 -256 8208 -160
rect 4864 -430 4870 -370
rect 4930 -377 5150 -370
rect 5462 -377 5513 -376
rect 7964 -377 7970 -370
rect 4930 -428 6540 -377
rect 7485 -428 7970 -377
rect 4930 -430 5150 -428
rect 5462 -494 5513 -428
rect 5462 -533 5468 -494
rect 5507 -533 5513 -494
rect 5462 -545 5513 -533
rect 5547 -493 5621 -487
rect 5547 -543 5559 -493
rect 5609 -543 5621 -493
rect 5547 -549 5621 -543
rect 7808 -494 7859 -428
rect 7964 -430 7970 -428
rect 8030 -377 8036 -370
rect 8030 -428 8040 -377
rect 8030 -430 8036 -428
rect 7808 -533 7814 -494
rect 7853 -533 7859 -494
rect 7808 -545 7859 -533
rect 7891 -493 7965 -487
rect 8610 -493 8770 -490
rect 7891 -543 7903 -493
rect 7953 -543 8770 -493
rect 7891 -549 7965 -543
rect 5314 -601 5320 -593
rect 5280 -651 5320 -601
rect 5314 -653 5320 -651
rect 5380 -601 5386 -593
rect 5559 -601 5609 -549
rect 8610 -550 8770 -543
rect 8830 -550 8836 -490
rect 5380 -651 5609 -601
rect 5380 -653 5386 -651
rect 5330 -800 8386 -704
rect 8482 -800 8488 -704
rect 3970 -1070 4410 -1010
rect 4470 -1070 4476 -1010
rect 5026 -1056 5032 -960
rect 5128 -1056 8165 -960
rect 4764 -1230 4770 -1170
rect 4830 -1177 5190 -1170
rect 8690 -1177 8890 -1170
rect 4830 -1228 6540 -1177
rect 7485 -1228 8890 -1177
rect 4830 -1230 5190 -1228
rect 5462 -1291 5513 -1228
rect 5462 -1330 5468 -1291
rect 5507 -1330 5513 -1291
rect 5462 -1342 5513 -1330
rect 5548 -1282 5622 -1276
rect 5548 -1332 5560 -1282
rect 5610 -1332 5622 -1282
rect 5548 -1338 5622 -1332
rect 7798 -1294 7849 -1228
rect 8690 -1230 8890 -1228
rect 8950 -1230 8956 -1170
rect 7798 -1333 7804 -1294
rect 7843 -1333 7849 -1294
rect 7891 -1277 7965 -1271
rect 7891 -1327 7903 -1277
rect 7953 -1290 8754 -1277
rect 7953 -1327 9010 -1290
rect 7891 -1333 7965 -1327
rect 2730 -1430 4290 -1370
rect 4350 -1430 4356 -1370
rect 4644 -1430 4650 -1370
rect 4710 -1390 5190 -1370
rect 5560 -1390 5610 -1338
rect 7798 -1345 7849 -1333
rect 8570 -1350 9010 -1327
rect 9070 -1350 9076 -1290
rect 4710 -1430 5610 -1390
rect 9180 -1410 9240 -1158
rect 2730 -1650 2790 -1430
rect 4935 -1440 5610 -1430
rect 8684 -1470 8690 -1410
rect 8750 -1470 9240 -1410
rect 5297 -1600 8398 -1504
rect 8494 -1600 8500 -1504
rect 11420 -1530 11480 -1158
rect 8804 -1590 8810 -1530
rect 8870 -1590 11480 -1530
rect 5046 -1856 5052 -1760
rect 5148 -1856 8183 -1760
rect 8924 -1798 8930 -1738
rect 8990 -1798 9350 -1738
rect 4524 -2030 4530 -1970
rect 4590 -1977 5270 -1970
rect 8684 -1977 8690 -1970
rect 4590 -2028 6540 -1977
rect 7485 -2028 8690 -1977
rect 4590 -2030 5270 -2028
rect 5460 -2092 5511 -2028
rect 5460 -2131 5466 -2092
rect 5505 -2131 5511 -2092
rect 5460 -2143 5511 -2131
rect 5548 -2082 5622 -2076
rect 5548 -2132 5560 -2082
rect 5610 -2132 5622 -2082
rect 5548 -2138 5622 -2132
rect 7807 -2091 7858 -2028
rect 8684 -2030 8690 -2028
rect 8750 -1977 8756 -1970
rect 8750 -2028 8760 -1977
rect 8750 -2030 8756 -2028
rect 7807 -2130 7813 -2091
rect 7852 -2130 7858 -2091
rect 4404 -2230 4410 -2170
rect 4470 -2190 5190 -2170
rect 5560 -2190 5610 -2138
rect 7807 -2142 7858 -2130
rect 7891 -2075 7965 -2069
rect 7891 -2125 7903 -2075
rect 7953 -2090 8800 -2075
rect 7953 -2125 8810 -2090
rect 7891 -2131 7965 -2125
rect 8690 -2150 8810 -2125
rect 8870 -2150 8876 -2090
rect 4470 -2230 5610 -2190
rect 5055 -2240 5610 -2230
rect 5312 -2400 8396 -2304
rect 8492 -2400 8498 -2304
rect 5040 -2655 5046 -2559
rect 5142 -2655 8154 -2559
rect 4070 -2970 4130 -2690
rect 4290 -2770 4350 -2764
rect 4350 -2777 5030 -2770
rect 8924 -2777 8930 -2770
rect 4350 -2828 6540 -2777
rect 7485 -2828 8930 -2777
rect 4350 -2830 5030 -2828
rect 4290 -2836 4350 -2830
rect 5458 -2892 5509 -2828
rect 5458 -2931 5464 -2892
rect 5503 -2931 5509 -2892
rect 5458 -2943 5509 -2931
rect 5548 -2882 5622 -2876
rect 5548 -2932 5560 -2882
rect 5610 -2932 5622 -2882
rect 5548 -2938 5622 -2932
rect 7802 -2892 7853 -2828
rect 8924 -2830 8930 -2828
rect 8990 -2830 8996 -2770
rect 7802 -2931 7808 -2892
rect 7847 -2931 7853 -2892
rect 4070 -2990 5070 -2970
rect 5560 -2990 5610 -2938
rect 7802 -2943 7853 -2931
rect 7891 -2883 7965 -2877
rect 7891 -2933 7903 -2883
rect 7953 -2890 8800 -2883
rect 7953 -2933 8730 -2890
rect 7891 -2939 7965 -2933
rect 8724 -2950 8730 -2933
rect 8790 -2933 8800 -2890
rect 8790 -2950 8796 -2933
rect 4070 -3030 5610 -2990
rect 4994 -3040 5610 -3030
rect 4850 -3090 4910 -3084
rect 2770 -3150 4850 -3090
rect 2770 -3350 2830 -3150
rect 4850 -3156 4910 -3150
rect 5344 -3200 8380 -3104
rect 8476 -3200 8482 -3104
rect 8724 -3162 8730 -3160
rect 8718 -3220 8730 -3162
rect 8790 -3162 8796 -3160
rect 11420 -3162 11480 -2850
rect 8790 -3220 11480 -3162
rect 8718 -3222 11480 -3220
rect 5056 -3456 5062 -3360
rect 5158 -3456 8208 -3360
rect 4844 -3630 4850 -3570
rect 4910 -3577 5070 -3570
rect 8770 -3577 9240 -3570
rect 4910 -3628 6540 -3577
rect 7485 -3628 9240 -3577
rect 4910 -3630 5070 -3628
rect 5451 -3693 5502 -3628
rect 5451 -3732 5457 -3693
rect 5496 -3732 5502 -3693
rect 5451 -3744 5502 -3732
rect 5548 -3678 5622 -3672
rect 5548 -3728 5560 -3678
rect 5610 -3728 5622 -3678
rect 5548 -3734 5622 -3728
rect 7802 -3694 7853 -3628
rect 8770 -3630 9240 -3628
rect 7802 -3733 7808 -3694
rect 7847 -3733 7853 -3694
rect 4070 -3786 5070 -3770
rect 5560 -3786 5610 -3734
rect 7802 -3745 7853 -3733
rect 7891 -3681 7965 -3675
rect 9014 -3680 9066 -3674
rect 7891 -3731 7903 -3681
rect 7953 -3731 9014 -3681
rect 7891 -3737 7965 -3731
rect 9014 -3738 9066 -3732
rect 4070 -3830 5610 -3786
rect 4994 -3836 5610 -3830
rect 5344 -4000 8370 -3904
rect 8466 -4000 8472 -3904
rect 5030 -4256 5036 -4160
rect 5132 -4256 8183 -4160
rect 8890 -4370 8950 -4364
rect 4204 -4430 4210 -4370
rect 4270 -4377 5110 -4370
rect 8730 -4377 8890 -4370
rect 4270 -4428 6540 -4377
rect 7485 -4428 8890 -4377
rect 4270 -4430 5110 -4428
rect 5460 -4492 5511 -4428
rect 5460 -4531 5466 -4492
rect 5505 -4531 5511 -4492
rect 5548 -4474 5622 -4468
rect 5548 -4524 5560 -4474
rect 5610 -4524 5622 -4474
rect 5548 -4530 5622 -4524
rect 7801 -4492 7852 -4428
rect 8730 -4430 8890 -4428
rect 8890 -4436 8950 -4430
rect 5460 -4543 5511 -4531
rect 4324 -4630 4330 -4570
rect 4390 -4582 5110 -4570
rect 5560 -4582 5610 -4530
rect 7801 -4531 7807 -4492
rect 7846 -4531 7852 -4492
rect 7801 -4543 7852 -4531
rect 7891 -4477 7965 -4471
rect 7891 -4527 7903 -4477
rect 7953 -4490 8825 -4477
rect 7953 -4527 8770 -4490
rect 7891 -4533 7965 -4527
rect 8764 -4550 8770 -4527
rect 8830 -4550 8836 -4490
rect 4390 -4630 5610 -4582
rect 4994 -4632 5610 -4630
rect 5297 -4800 8388 -4704
rect 8484 -4800 8490 -4704
rect 9008 -4730 9338 -4728
rect 9002 -4790 9010 -4730
rect 9070 -4788 9338 -4730
rect 9070 -4790 9096 -4788
rect 9002 -4796 9096 -4790
rect 2730 -4870 4210 -4810
rect 4270 -4870 4276 -4810
rect 9278 -4866 9338 -4788
rect 11420 -4866 11480 -4558
rect 2730 -5050 2790 -4870
rect 8874 -4890 8968 -4882
rect 8874 -4948 8890 -4890
rect 8878 -4950 8890 -4948
rect 8950 -4896 8968 -4890
rect 8950 -4950 9240 -4896
rect 9278 -4926 11480 -4866
rect 8878 -4956 9240 -4950
rect 4070 -5050 4330 -4990
rect 4390 -5050 4396 -4990
rect 5030 -5056 5036 -4960
rect 5132 -5056 8172 -4960
rect 8770 -5010 8830 -5004
rect 8830 -5070 9010 -5010
rect 9070 -5070 9076 -5010
rect 8770 -5076 8830 -5070
rect 4244 -5230 4250 -5170
rect 4310 -5177 5070 -5170
rect 8370 -5177 8890 -5170
rect 4310 -5228 6540 -5177
rect 7485 -5228 8890 -5177
rect 4310 -5230 5070 -5228
rect 5458 -5291 5509 -5228
rect 5458 -5330 5464 -5291
rect 5503 -5330 5509 -5291
rect 5458 -5342 5509 -5330
rect 5548 -5276 5622 -5270
rect 5548 -5326 5560 -5276
rect 5610 -5326 5622 -5276
rect 5548 -5332 5622 -5326
rect 7796 -5290 7847 -5228
rect 8370 -5230 8890 -5228
rect 8950 -5230 8956 -5170
rect 9180 -5208 9240 -4956
rect 7796 -5329 7802 -5290
rect 7841 -5329 7847 -5290
rect 4364 -5430 4370 -5370
rect 4430 -5384 5150 -5370
rect 5560 -5384 5610 -5332
rect 7796 -5341 7847 -5329
rect 7891 -5277 7965 -5271
rect 7891 -5327 7903 -5277
rect 7953 -5290 8560 -5277
rect 7953 -5327 8770 -5290
rect 7891 -5333 7965 -5327
rect 8410 -5350 8770 -5327
rect 8830 -5350 8836 -5290
rect 4430 -5430 5610 -5384
rect 4994 -5434 5610 -5430
rect 5337 -5600 8370 -5504
rect 8466 -5600 8472 -5504
rect 5026 -5856 5032 -5760
rect 5128 -5856 8201 -5760
rect 4484 -6030 4490 -5970
rect 4550 -5977 5070 -5970
rect 8090 -5977 8130 -5970
rect 4550 -6028 6540 -5977
rect 7485 -6028 8130 -5977
rect 4550 -6030 5070 -6028
rect 5457 -6093 5508 -6028
rect 5457 -6132 5463 -6093
rect 5502 -6132 5508 -6093
rect 5548 -6070 5622 -6064
rect 5548 -6120 5560 -6070
rect 5610 -6090 5622 -6070
rect 5548 -6126 5570 -6120
rect 5457 -6144 5508 -6132
rect 5560 -6150 5570 -6126
rect 5630 -6150 5636 -6090
rect 7801 -6095 7852 -6028
rect 8090 -6030 8130 -6028
rect 8190 -5977 8196 -5970
rect 8190 -6028 8200 -5977
rect 8190 -6030 8196 -6028
rect 7801 -6134 7807 -6095
rect 7846 -6134 7852 -6095
rect 7801 -6146 7852 -6134
rect 7891 -6087 7965 -6081
rect 7891 -6137 7903 -6087
rect 7953 -6090 8560 -6087
rect 8650 -6090 8710 -6084
rect 7953 -6137 8650 -6090
rect 7891 -6143 7965 -6137
rect 8410 -6150 8650 -6137
rect 5560 -6178 5610 -6150
rect 8650 -6156 8710 -6150
rect 5305 -6399 8394 -6303
rect 8490 -6399 8496 -6303
rect 2770 -6470 4250 -6410
rect 4310 -6470 4316 -6410
rect 2770 -6750 2830 -6470
rect 11420 -6562 11480 -6250
rect 9004 -6622 9010 -6562
rect 9070 -6622 11480 -6562
rect 3970 -6750 4370 -6690
rect 4430 -6750 4436 -6690
rect 8884 -6898 8890 -6838
rect 8950 -6898 9350 -6838
rect 5026 -7044 5032 -6948
rect 5128 -7044 7956 -6948
rect 6622 -7200 6706 -7194
rect 6065 -7260 6125 -7254
rect 6063 -7316 6065 -7264
rect 6195 -7260 6255 -7254
rect 6125 -7316 6127 -7264
rect 6193 -7316 6195 -7264
rect 6345 -7260 6405 -7254
rect 6065 -7326 6125 -7320
rect 6255 -7316 6257 -7264
rect 6343 -7316 6345 -7264
rect 6475 -7260 6535 -7254
rect 6195 -7326 6255 -7320
rect 6405 -7316 6407 -7264
rect 6473 -7316 6475 -7264
rect 6622 -7260 6634 -7200
rect 6694 -7260 6706 -7200
rect 7522 -7200 7606 -7194
rect 6345 -7326 6405 -7320
rect 6535 -7316 6537 -7264
rect 6622 -7266 6706 -7260
rect 6953 -7264 7013 -7258
rect 6951 -7320 6953 -7268
rect 7083 -7264 7143 -7258
rect 6475 -7326 6535 -7320
rect 6622 -7328 6706 -7322
rect 6622 -7388 6634 -7328
rect 6694 -7388 6706 -7328
rect 7013 -7320 7015 -7268
rect 7081 -7320 7083 -7268
rect 7233 -7264 7293 -7258
rect 6953 -7330 7013 -7324
rect 7143 -7320 7145 -7268
rect 7231 -7320 7233 -7268
rect 7363 -7264 7423 -7258
rect 7083 -7330 7143 -7324
rect 7293 -7320 7295 -7268
rect 7361 -7320 7363 -7268
rect 7522 -7260 7534 -7200
rect 7594 -7260 7606 -7200
rect 7522 -7266 7606 -7260
rect 7233 -7330 7293 -7324
rect 7423 -7320 7425 -7268
rect 7363 -7330 7423 -7324
rect 7522 -7328 7606 -7322
rect 6622 -7394 6706 -7388
rect 7522 -7388 7534 -7328
rect 7594 -7388 7606 -7328
rect 7522 -7394 7606 -7388
rect 5682 -7582 8372 -7486
rect 8468 -7582 8474 -7486
rect 8768 -8170 9368 -8164
rect 4490 -8210 4550 -8204
rect 8764 -8230 8770 -8170
rect 8830 -8224 9368 -8170
rect 8830 -8230 8848 -8224
rect 8764 -8236 8848 -8230
rect 4490 -8598 4550 -8270
rect 9308 -8264 9368 -8224
rect 11420 -8264 11480 -7930
rect 9308 -8324 11480 -8264
rect 8650 -8330 8710 -8324
rect 8130 -8370 8190 -8364
rect 5564 -8430 5570 -8370
rect 5630 -8430 5636 -8370
rect 8710 -8390 9280 -8330
rect 8650 -8396 8710 -8390
rect 5570 -8598 5630 -8430
rect 8130 -8598 8190 -8430
rect 9220 -8598 9280 -8390
<< via1 >>
rect 5320 1996 5380 2060
rect 4768 1868 4828 1928
rect 4870 1870 4930 1930
rect 7970 1806 8030 1866
rect 8770 1824 8830 1884
rect 8890 1602 8950 1662
rect 5042 984 5138 1080
rect 5876 814 5946 824
rect 5876 764 5946 814
rect 7504 760 7564 820
rect 6036 744 6096 754
rect 6036 704 6046 744
rect 6046 704 6086 744
rect 6086 704 6096 744
rect 4650 630 4710 690
rect 5876 634 5946 694
rect 6036 694 6096 704
rect 6166 744 6226 754
rect 6166 704 6176 744
rect 6176 704 6216 744
rect 6216 704 6226 744
rect 6166 694 6226 704
rect 6316 744 6376 754
rect 6316 704 6326 744
rect 6326 704 6366 744
rect 6366 704 6376 744
rect 6316 694 6376 704
rect 6446 744 6506 754
rect 6446 704 6456 744
rect 6456 704 6496 744
rect 6496 704 6506 744
rect 6446 694 6506 704
rect 6926 744 6986 754
rect 6926 704 6936 744
rect 6936 704 6976 744
rect 6976 704 6986 744
rect 6926 694 6986 704
rect 7056 744 7116 754
rect 7056 704 7066 744
rect 7066 704 7106 744
rect 7106 704 7116 744
rect 7056 694 7116 704
rect 7206 744 7266 754
rect 7206 704 7216 744
rect 7216 704 7256 744
rect 7256 704 7266 744
rect 7206 694 7266 704
rect 7336 744 7396 754
rect 7336 704 7346 744
rect 7346 704 7386 744
rect 7386 704 7396 744
rect 7336 694 7396 704
rect 7503 631 7572 700
rect 8416 440 8512 536
rect 4530 250 4590 310
rect 9010 136 9070 196
rect 5062 -256 5158 -160
rect 4870 -430 4930 -370
rect 7970 -430 8030 -370
rect 5320 -653 5380 -593
rect 8770 -550 8830 -490
rect 8386 -800 8482 -704
rect 4410 -1070 4470 -1010
rect 5032 -1056 5128 -960
rect 4770 -1230 4830 -1170
rect 8890 -1230 8950 -1170
rect 4290 -1430 4350 -1370
rect 4650 -1430 4710 -1370
rect 9010 -1350 9070 -1290
rect 8690 -1470 8750 -1410
rect 8398 -1600 8494 -1504
rect 8810 -1590 8870 -1530
rect 5052 -1856 5148 -1760
rect 8930 -1798 8990 -1738
rect 4530 -2030 4590 -1970
rect 8690 -2030 8750 -1970
rect 4410 -2230 4470 -2170
rect 8810 -2150 8870 -2090
rect 8396 -2400 8492 -2304
rect 5046 -2655 5142 -2559
rect 4290 -2830 4350 -2770
rect 8930 -2830 8990 -2770
rect 8730 -2950 8790 -2890
rect 4850 -3150 4910 -3090
rect 8380 -3200 8476 -3104
rect 8730 -3220 8790 -3160
rect 5062 -3456 5158 -3360
rect 4850 -3630 4910 -3570
rect 9014 -3732 9066 -3680
rect 8370 -4000 8466 -3904
rect 5036 -4256 5132 -4160
rect 4210 -4430 4270 -4370
rect 8890 -4430 8950 -4370
rect 4330 -4630 4390 -4570
rect 8770 -4550 8830 -4490
rect 8388 -4800 8484 -4704
rect 9010 -4790 9070 -4730
rect 4210 -4870 4270 -4810
rect 8890 -4950 8950 -4890
rect 4330 -5050 4390 -4990
rect 5036 -5056 5132 -4960
rect 8770 -5070 8830 -5010
rect 9010 -5070 9070 -5010
rect 4250 -5230 4310 -5170
rect 8890 -5230 8950 -5170
rect 4370 -5430 4430 -5370
rect 8770 -5350 8830 -5290
rect 8370 -5600 8466 -5504
rect 5032 -5856 5128 -5760
rect 4490 -6030 4550 -5970
rect 5570 -6120 5610 -6090
rect 5610 -6120 5630 -6090
rect 5570 -6150 5630 -6120
rect 8130 -6030 8190 -5970
rect 8650 -6150 8710 -6090
rect 8394 -6399 8490 -6303
rect 4250 -6470 4310 -6410
rect 9010 -6622 9070 -6562
rect 4370 -6750 4430 -6690
rect 8890 -6898 8950 -6838
rect 5032 -7044 5128 -6948
rect 6065 -7270 6125 -7260
rect 6065 -7310 6075 -7270
rect 6075 -7310 6115 -7270
rect 6115 -7310 6125 -7270
rect 6065 -7320 6125 -7310
rect 6195 -7270 6255 -7260
rect 6195 -7310 6205 -7270
rect 6205 -7310 6245 -7270
rect 6245 -7310 6255 -7270
rect 6195 -7320 6255 -7310
rect 6345 -7270 6405 -7260
rect 6345 -7310 6355 -7270
rect 6355 -7310 6395 -7270
rect 6395 -7310 6405 -7270
rect 6345 -7320 6405 -7310
rect 6475 -7270 6535 -7260
rect 6634 -7260 6694 -7200
rect 6475 -7310 6485 -7270
rect 6485 -7310 6525 -7270
rect 6525 -7310 6535 -7270
rect 6475 -7320 6535 -7310
rect 6953 -7274 7013 -7264
rect 6953 -7314 6963 -7274
rect 6963 -7314 7003 -7274
rect 7003 -7314 7013 -7274
rect 6634 -7388 6694 -7328
rect 6953 -7324 7013 -7314
rect 7083 -7274 7143 -7264
rect 7083 -7314 7093 -7274
rect 7093 -7314 7133 -7274
rect 7133 -7314 7143 -7274
rect 7083 -7324 7143 -7314
rect 7233 -7274 7293 -7264
rect 7233 -7314 7243 -7274
rect 7243 -7314 7283 -7274
rect 7283 -7314 7293 -7274
rect 7233 -7324 7293 -7314
rect 7363 -7274 7423 -7264
rect 7534 -7260 7594 -7200
rect 7363 -7314 7373 -7274
rect 7373 -7314 7413 -7274
rect 7413 -7314 7423 -7274
rect 7363 -7324 7423 -7314
rect 7534 -7388 7594 -7328
rect 8372 -7582 8468 -7486
rect 4490 -8270 4550 -8210
rect 8770 -8230 8830 -8170
rect 5570 -8430 5630 -8370
rect 8130 -8430 8190 -8370
rect 8650 -8390 8710 -8330
<< metal2 >>
rect 12953 3254 13207 3263
rect 184 3000 193 3254
rect 447 3000 5407 3254
rect 8993 3000 12953 3254
rect 12953 2991 13207 3000
rect -327 2328 5427 2582
rect 8973 2328 13727 2582
rect 5314 1996 5320 2060
rect 5380 1996 5386 2060
rect 4870 1930 4930 1936
rect 4762 1868 4768 1928
rect 4828 1868 4834 1928
rect 4768 1864 4830 1868
rect 184 1420 193 1674
rect 447 1420 3047 1674
rect -327 748 3027 1002
rect 4650 690 4710 696
rect 4524 250 4530 310
rect 4590 250 4596 310
rect 184 -280 193 -26
rect 447 -280 3047 -26
rect -327 -952 3027 -698
rect 4410 -1010 4470 -1004
rect 4290 -1370 4350 -1364
rect 184 -1980 193 -1726
rect 447 -1980 3047 -1726
rect -327 -2652 3027 -2398
rect 4290 -2770 4350 -1430
rect 4410 -2170 4470 -1070
rect 4530 -1970 4590 250
rect 4650 -1370 4710 630
rect 4770 -1170 4830 1864
rect 4870 -370 4930 1870
rect 5042 1080 5138 1090
rect 5042 974 5138 984
rect 5062 -160 5158 -150
rect 5062 -266 5158 -256
rect 4870 -436 4930 -430
rect 5320 -593 5380 1996
rect 8770 1884 8830 1890
rect 7970 1866 8030 1872
rect 5876 824 5946 834
rect 5876 700 5946 764
rect 7504 820 7564 830
rect 5870 694 5946 700
rect 5996 694 6036 754
rect 6096 694 6166 754
rect 6226 694 6316 754
rect 6376 694 6446 754
rect 6506 694 6566 754
rect 6886 694 6926 754
rect 6986 694 7056 754
rect 7116 694 7206 754
rect 7266 694 7336 754
rect 7396 694 7456 754
rect 7504 710 7564 760
rect 7503 700 7572 710
rect 5870 684 5876 694
rect 5866 634 5876 684
rect 5866 624 5946 634
rect 5870 458 5930 624
rect 6166 602 6226 694
rect 7040 604 7100 694
rect 7503 621 7572 631
rect 6159 546 6168 602
rect 6224 546 6233 602
rect 7033 548 7042 604
rect 7098 548 7107 604
rect 7040 546 7100 548
rect 6166 544 6226 546
rect 5863 402 5872 458
rect 5928 402 5937 458
rect 5870 400 5930 402
rect 7504 372 7564 621
rect 7504 316 7506 372
rect 7562 316 7564 372
rect 7504 314 7564 316
rect 7506 307 7562 314
rect 6130 208 7170 210
rect 6123 152 6132 208
rect 6188 152 7170 208
rect 6130 150 7170 152
rect 7230 150 7239 210
rect 6000 118 7040 120
rect 5993 62 6002 118
rect 6058 62 7040 118
rect 6000 60 7040 62
rect 7100 60 7109 120
rect 5870 28 6910 30
rect 5863 -28 5872 28
rect 5928 -28 6910 28
rect 5870 -30 6910 -28
rect 6970 -30 6979 30
rect 5740 -62 6780 -60
rect 5733 -118 5742 -62
rect 5798 -118 6780 -62
rect 5740 -120 6780 -118
rect 6840 -120 6849 -60
rect 7970 -370 8030 1806
rect 8416 536 8512 546
rect 8416 430 8512 440
rect 7970 -436 8030 -430
rect 6392 -482 6448 -475
rect 6034 -484 6190 -482
rect 6308 -484 6450 -482
rect 6780 -484 6910 -482
rect 5863 -546 5872 -490
rect 5928 -546 5937 -490
rect 6034 -540 6132 -484
rect 6188 -540 6197 -484
rect 6308 -540 6392 -484
rect 6448 -540 6450 -484
rect 6034 -542 6190 -540
rect 6308 -542 6450 -540
rect 6643 -542 6652 -486
rect 6708 -542 6717 -486
rect 6773 -540 6782 -484
rect 6838 -540 6910 -484
rect 6780 -542 6910 -540
rect 6392 -549 6448 -542
rect 7033 -552 7042 -496
rect 7098 -552 7107 -496
rect 7293 -546 7302 -490
rect 7358 -546 7367 -490
rect 7620 -564 7680 -482
rect 8770 -490 8830 1824
rect 8770 -556 8830 -550
rect 8890 1662 8950 1668
rect 7560 -566 7680 -564
rect 7553 -622 7562 -566
rect 7618 -622 7680 -566
rect 7560 -624 7680 -622
rect 5320 -659 5380 -653
rect 8386 -704 8482 -694
rect 8386 -810 8482 -800
rect 5032 -960 5128 -950
rect 5032 -1066 5128 -1056
rect 4770 -1236 4830 -1230
rect 8890 -1170 8950 1602
rect 11273 1272 12953 1526
rect 13207 1272 13216 1526
rect 11273 600 13727 854
rect 9010 196 9070 208
rect 9004 136 9010 196
rect 9070 136 9076 196
rect 8890 -1236 8950 -1230
rect 6306 -1288 6450 -1286
rect 6652 -1288 6708 -1279
rect 6038 -1290 6190 -1288
rect 5740 -1292 5912 -1290
rect 5733 -1348 5742 -1292
rect 5798 -1348 5912 -1292
rect 6038 -1346 6132 -1290
rect 6188 -1346 6197 -1290
rect 6306 -1344 6392 -1288
rect 6448 -1344 6457 -1288
rect 6306 -1346 6450 -1344
rect 6038 -1348 6190 -1346
rect 5740 -1350 5912 -1348
rect 6652 -1353 6708 -1344
rect 6848 -1292 6970 -1290
rect 6848 -1348 6912 -1292
rect 6968 -1348 6977 -1292
rect 7033 -1342 7042 -1286
rect 7098 -1342 7107 -1286
rect 9010 -1290 9070 136
rect 11233 -428 12953 -174
rect 13207 -428 13216 -174
rect 11273 -1100 13727 -846
rect 7293 -1346 7302 -1290
rect 7358 -1346 7367 -1290
rect 6848 -1350 6970 -1348
rect 7614 -1382 7674 -1290
rect 9010 -1356 9070 -1350
rect 7560 -1384 7674 -1382
rect 4650 -1436 4710 -1430
rect 7553 -1440 7562 -1384
rect 7618 -1440 7674 -1384
rect 7560 -1442 7674 -1440
rect 8690 -1410 8750 -1404
rect 8398 -1504 8494 -1494
rect 8398 -1610 8494 -1600
rect 5052 -1760 5148 -1750
rect 5052 -1866 5148 -1856
rect 4530 -2036 4590 -2030
rect 8690 -1970 8750 -1470
rect 8690 -2036 8750 -2030
rect 8810 -1530 8870 -1524
rect 5863 -2142 5872 -2086
rect 5928 -2142 5937 -2086
rect 6324 -2088 6450 -2086
rect 5993 -2148 6002 -2092
rect 6058 -2148 6067 -2092
rect 6324 -2144 6392 -2088
rect 6448 -2144 6457 -2088
rect 6643 -2138 6652 -2082
rect 6708 -2138 6717 -2082
rect 6780 -2092 6906 -2090
rect 6324 -2146 6450 -2144
rect 6773 -2148 6782 -2092
rect 6838 -2148 6906 -2092
rect 6780 -2150 6906 -2148
rect 7032 -2094 7230 -2092
rect 7032 -2150 7172 -2094
rect 7228 -2150 7237 -2094
rect 7293 -2144 7302 -2088
rect 7358 -2144 7367 -2088
rect 8810 -2090 8870 -1590
rect 7032 -2152 7230 -2150
rect 7614 -2166 7674 -2100
rect 8810 -2156 8870 -2150
rect 8930 -1738 8990 -1732
rect 7560 -2168 7674 -2166
rect 7553 -2224 7562 -2168
rect 7618 -2224 7674 -2168
rect 7560 -2226 7674 -2224
rect 4410 -2236 4470 -2230
rect 8396 -2304 8492 -2294
rect 8396 -2410 8492 -2400
rect 5046 -2559 5142 -2549
rect 5046 -2665 5142 -2655
rect 8930 -2770 8990 -1798
rect 11233 -2128 12953 -1874
rect 13207 -2128 13216 -1874
rect 4284 -2830 4290 -2770
rect 4350 -2830 4356 -2770
rect 11273 -2800 13727 -2546
rect 8930 -2836 8990 -2830
rect 5740 -2884 5904 -2882
rect 5733 -2940 5742 -2884
rect 5798 -2940 5904 -2884
rect 5740 -2942 5904 -2940
rect 5993 -2942 6002 -2886
rect 6058 -2942 6067 -2886
rect 6320 -2890 6450 -2888
rect 6320 -2946 6392 -2890
rect 6448 -2946 6457 -2890
rect 6643 -2944 6652 -2888
rect 6708 -2944 6717 -2888
rect 6850 -2892 6970 -2890
rect 6320 -2948 6450 -2946
rect 6850 -2948 6912 -2892
rect 6968 -2948 6977 -2892
rect 7026 -2898 7230 -2896
rect 6850 -2950 6970 -2948
rect 7026 -2954 7172 -2898
rect 7228 -2954 7237 -2898
rect 7293 -2940 7302 -2884
rect 7358 -2940 7367 -2884
rect 7026 -2956 7230 -2954
rect 7620 -2980 7680 -2888
rect 7560 -2982 7680 -2980
rect 7553 -3038 7562 -2982
rect 7618 -3038 7680 -2982
rect 7560 -3040 7680 -3038
rect 8730 -2890 8790 -2884
rect 4844 -3150 4850 -3090
rect 4910 -3150 4916 -3090
rect 8380 -3104 8476 -3094
rect 184 -3680 193 -3426
rect 447 -3680 3007 -3426
rect 4850 -3570 4910 -3150
rect 8380 -3210 8476 -3200
rect 8730 -3160 8790 -2950
rect 8730 -3226 8790 -3220
rect 5062 -3360 5158 -3350
rect 5062 -3466 5158 -3456
rect 4850 -3636 4910 -3630
rect 9010 -3680 9070 -3650
rect 5863 -3740 5872 -3684
rect 5928 -3740 5937 -3684
rect 6054 -3688 6190 -3686
rect 6054 -3744 6132 -3688
rect 6188 -3744 6197 -3688
rect 6253 -3740 6262 -3684
rect 6318 -3740 6327 -3684
rect 6054 -3746 6190 -3744
rect 6643 -3746 6652 -3690
rect 6708 -3746 6717 -3690
rect 6780 -3694 6906 -3692
rect 6773 -3750 6782 -3694
rect 6838 -3750 6906 -3694
rect 6780 -3752 6906 -3750
rect 7033 -3754 7042 -3698
rect 7098 -3754 7107 -3698
rect 7304 -3770 7364 -3694
rect 7432 -3770 7488 -3763
rect 7304 -3772 7490 -3770
rect 7304 -3828 7432 -3772
rect 7488 -3828 7490 -3772
rect 7618 -3774 7678 -3682
rect 9008 -3732 9014 -3680
rect 9066 -3732 9072 -3680
rect 7560 -3776 7678 -3774
rect 7304 -3830 7490 -3828
rect 7432 -3837 7488 -3830
rect 7553 -3832 7562 -3776
rect 7618 -3832 7678 -3776
rect 7560 -3834 7678 -3832
rect 8370 -3904 8466 -3894
rect 8370 -4010 8466 -4000
rect -327 -4352 3027 -4098
rect 5036 -4160 5132 -4150
rect 5036 -4266 5132 -4256
rect 4210 -4370 4270 -4364
rect 8884 -4430 8890 -4370
rect 8950 -4430 8956 -4370
rect 4210 -4810 4270 -4430
rect 6052 -4488 6190 -4486
rect 5740 -4496 5916 -4494
rect 5733 -4552 5742 -4496
rect 5798 -4552 5916 -4496
rect 6052 -4544 6132 -4488
rect 6188 -4544 6197 -4488
rect 6052 -4546 6190 -4544
rect 6253 -4548 6262 -4492
rect 6318 -4548 6327 -4492
rect 6643 -4542 6652 -4486
rect 6708 -4542 6717 -4486
rect 6858 -4488 6970 -4486
rect 6858 -4544 6912 -4488
rect 6968 -4544 6977 -4488
rect 7033 -4542 7042 -4486
rect 7098 -4542 7107 -4486
rect 6858 -4546 6970 -4544
rect 5740 -4554 5916 -4552
rect 4210 -4876 4270 -4870
rect 4330 -4570 4390 -4564
rect 4330 -4990 4390 -4630
rect 7298 -4572 7358 -4492
rect 7432 -4572 7488 -4565
rect 7616 -4570 7676 -4486
rect 7560 -4572 7676 -4570
rect 7298 -4574 7490 -4572
rect 7298 -4630 7432 -4574
rect 7488 -4630 7490 -4574
rect 7553 -4628 7562 -4572
rect 7618 -4628 7676 -4572
rect 7560 -4630 7676 -4628
rect 8770 -4490 8830 -4484
rect 7298 -4632 7490 -4630
rect 7432 -4639 7488 -4632
rect 8388 -4704 8484 -4694
rect 8388 -4810 8484 -4800
rect 4330 -5056 4390 -5050
rect 5036 -4960 5132 -4950
rect 8770 -5010 8830 -4550
rect 8890 -4890 8950 -4430
rect 9010 -4730 9070 -3732
rect 11273 -3828 12953 -3574
rect 13207 -3828 13216 -3574
rect 11273 -4500 13727 -4246
rect 9010 -4796 9070 -4790
rect 8890 -4956 8950 -4950
rect 9010 -5010 9070 -5004
rect 5036 -5066 5132 -5056
rect 8764 -5070 8770 -5010
rect 8830 -5070 8836 -5010
rect 184 -5380 193 -5126
rect 447 -5380 3047 -5126
rect 4250 -5170 4310 -5164
rect -327 -6052 3027 -5798
rect 4250 -6410 4310 -5230
rect 8890 -5170 8950 -5164
rect 5863 -5346 5872 -5290
rect 5928 -5346 5937 -5290
rect 6780 -5292 6902 -5290
rect 5993 -5348 6002 -5292
rect 6058 -5348 6067 -5292
rect 6253 -5350 6262 -5294
rect 6318 -5350 6327 -5294
rect 6643 -5348 6652 -5292
rect 6708 -5348 6717 -5292
rect 6773 -5348 6782 -5292
rect 6838 -5348 6902 -5292
rect 6780 -5350 6902 -5348
rect 7032 -5296 7230 -5294
rect 7032 -5352 7172 -5296
rect 7228 -5352 7237 -5296
rect 7032 -5354 7230 -5352
rect 4250 -6476 4310 -6470
rect 4370 -5370 4430 -5364
rect 4370 -6690 4430 -5430
rect 7314 -5382 7374 -5296
rect 7620 -5380 7680 -5288
rect 7560 -5382 7680 -5380
rect 7314 -5384 7490 -5382
rect 7314 -5440 7432 -5384
rect 7488 -5440 7497 -5384
rect 7553 -5438 7562 -5382
rect 7618 -5438 7680 -5382
rect 7560 -5440 7680 -5438
rect 8770 -5290 8830 -5284
rect 7314 -5442 7490 -5440
rect 8370 -5504 8466 -5494
rect 8370 -5610 8466 -5600
rect 5032 -5760 5128 -5750
rect 5032 -5866 5128 -5856
rect 4370 -6756 4430 -6750
rect 4490 -5970 4550 -5964
rect 184 -7080 193 -6826
rect 447 -7080 3047 -6826
rect -327 -7752 3027 -7498
rect 4490 -8210 4550 -6030
rect 8130 -5970 8190 -5964
rect 7022 -6082 7230 -6080
rect 5570 -6090 5630 -6084
rect 5740 -6102 5908 -6100
rect 5032 -6948 5128 -6938
rect 5032 -7054 5128 -7044
rect 4484 -8270 4490 -8210
rect 4550 -8270 4556 -8210
rect 5570 -8370 5630 -6150
rect 5733 -6158 5742 -6102
rect 5798 -6158 5908 -6102
rect 5993 -6146 6002 -6090
rect 6058 -6146 6067 -6090
rect 6253 -6146 6262 -6090
rect 6318 -6146 6327 -6090
rect 6643 -6142 6652 -6086
rect 6708 -6142 6717 -6086
rect 6838 -6090 6970 -6088
rect 6838 -6146 6912 -6090
rect 6968 -6146 6977 -6090
rect 7022 -6138 7172 -6082
rect 7228 -6138 7237 -6082
rect 7022 -6140 7230 -6138
rect 6838 -6148 6970 -6146
rect 5740 -6160 5908 -6158
rect 7304 -6176 7364 -6090
rect 7304 -6178 7490 -6176
rect 7304 -6234 7432 -6178
rect 7488 -6234 7497 -6178
rect 7618 -6180 7678 -6094
rect 7560 -6182 7678 -6180
rect 7304 -6236 7490 -6234
rect 7553 -6238 7562 -6182
rect 7618 -6238 7678 -6182
rect 7560 -6240 7678 -6238
rect 6260 -6452 7300 -6450
rect 6253 -6508 6262 -6452
rect 6318 -6508 7300 -6452
rect 6260 -6510 7300 -6508
rect 7360 -6510 7369 -6450
rect 6390 -6542 7430 -6540
rect 6383 -6598 6392 -6542
rect 6448 -6598 7430 -6542
rect 6390 -6600 7430 -6598
rect 7490 -6600 7499 -6540
rect 6520 -6632 7560 -6630
rect 6513 -6688 6522 -6632
rect 6578 -6688 7560 -6632
rect 6520 -6690 7560 -6688
rect 7620 -6690 7629 -6630
rect 6650 -6722 7690 -6720
rect 6643 -6778 6652 -6722
rect 6708 -6778 7690 -6722
rect 6650 -6780 7690 -6778
rect 7750 -6780 7759 -6720
rect 7158 -7002 7214 -6995
rect 7156 -7004 7216 -7002
rect 6634 -7052 6694 -7050
rect 6260 -7058 6320 -7056
rect 6253 -7114 6262 -7058
rect 6318 -7114 6327 -7058
rect 6627 -7108 6636 -7052
rect 6692 -7108 6701 -7052
rect 7156 -7060 7158 -7004
rect 7214 -7060 7216 -7004
rect 6260 -7260 6320 -7114
rect 6634 -7200 6694 -7108
rect 6025 -7320 6065 -7260
rect 6125 -7320 6195 -7260
rect 6255 -7320 6345 -7260
rect 6405 -7320 6475 -7260
rect 6535 -7320 6595 -7260
rect 6634 -7328 6694 -7260
rect 7156 -7264 7216 -7060
rect 7534 -7198 7594 -7194
rect 7534 -7200 7750 -7198
rect 7594 -7256 7692 -7200
rect 7748 -7256 7757 -7200
rect 7594 -7258 7750 -7256
rect 6913 -7324 6953 -7264
rect 7013 -7324 7083 -7264
rect 7143 -7324 7233 -7264
rect 7293 -7324 7363 -7264
rect 7423 -7324 7483 -7264
rect 6634 -7394 6694 -7388
rect 7534 -7328 7594 -7260
rect 7534 -7394 7594 -7388
rect 8130 -8370 8190 -6030
rect 8644 -6150 8650 -6090
rect 8710 -6150 8716 -6090
rect 8394 -6303 8490 -6293
rect 8394 -6409 8490 -6399
rect 8372 -7486 8468 -7476
rect 8372 -7592 8468 -7582
rect 8650 -8330 8710 -6150
rect 8770 -8170 8830 -5350
rect 8890 -6838 8950 -5230
rect 9010 -6562 9070 -5070
rect 11273 -5528 12953 -5274
rect 13207 -5528 13216 -5274
rect 11273 -6200 13727 -5946
rect 9010 -6628 9070 -6622
rect 8890 -6904 8950 -6898
rect 11273 -7228 12953 -6974
rect 13207 -7228 13216 -6974
rect 11273 -7900 13727 -7646
rect 8770 -8236 8830 -8230
rect 8124 -8430 8130 -8370
rect 8190 -8430 8196 -8370
rect 8644 -8390 8650 -8330
rect 8710 -8390 8716 -8330
rect 5570 -8436 5630 -8430
rect 184 -8928 193 -8674
rect 447 -8928 5527 -8674
rect 9033 -8928 12953 -8674
rect 13207 -8928 13216 -8674
rect -327 -9600 5527 -9346
rect 9073 -9600 13727 -9346
<< via2 >>
rect 193 3000 447 3254
rect 12953 3000 13207 3254
rect 193 1420 447 1674
rect 193 -280 447 -26
rect 193 -1980 447 -1726
rect 5042 984 5138 1080
rect 5062 -256 5158 -160
rect 6168 546 6224 602
rect 7042 548 7098 604
rect 5872 402 5928 458
rect 7506 316 7562 372
rect 6132 152 6188 208
rect 7170 150 7230 210
rect 6002 62 6058 118
rect 7040 60 7100 120
rect 5872 -28 5928 28
rect 6910 -30 6970 30
rect 5742 -118 5798 -62
rect 6780 -120 6840 -60
rect 8416 440 8512 536
rect 5872 -546 5928 -490
rect 6132 -540 6188 -484
rect 6392 -540 6448 -484
rect 6652 -542 6708 -486
rect 6782 -540 6838 -484
rect 7042 -552 7098 -496
rect 7302 -546 7358 -490
rect 7562 -622 7618 -566
rect 8386 -800 8482 -704
rect 5032 -1056 5128 -960
rect 12953 1272 13207 1526
rect 5742 -1348 5798 -1292
rect 6132 -1346 6188 -1290
rect 6392 -1344 6448 -1288
rect 6652 -1344 6708 -1288
rect 6912 -1348 6968 -1292
rect 7042 -1342 7098 -1286
rect 12953 -428 13207 -174
rect 7302 -1346 7358 -1290
rect 7562 -1440 7618 -1384
rect 8398 -1600 8494 -1504
rect 5052 -1856 5148 -1760
rect 5872 -2142 5928 -2086
rect 6002 -2148 6058 -2092
rect 6392 -2144 6448 -2088
rect 6652 -2138 6708 -2082
rect 6782 -2148 6838 -2092
rect 7172 -2150 7228 -2094
rect 7302 -2144 7358 -2088
rect 7562 -2224 7618 -2168
rect 8396 -2400 8492 -2304
rect 5046 -2655 5142 -2559
rect 12953 -2128 13207 -1874
rect 5742 -2940 5798 -2884
rect 6002 -2942 6058 -2886
rect 6392 -2946 6448 -2890
rect 6652 -2944 6708 -2888
rect 6912 -2948 6968 -2892
rect 7172 -2954 7228 -2898
rect 7302 -2940 7358 -2884
rect 7562 -3038 7618 -2982
rect 193 -3680 447 -3426
rect 8380 -3200 8476 -3104
rect 5062 -3456 5158 -3360
rect 5872 -3740 5928 -3684
rect 6132 -3744 6188 -3688
rect 6262 -3740 6318 -3684
rect 6652 -3746 6708 -3690
rect 6782 -3750 6838 -3694
rect 7042 -3754 7098 -3698
rect 7432 -3828 7488 -3772
rect 7562 -3832 7618 -3776
rect 8370 -4000 8466 -3904
rect 5036 -4256 5132 -4160
rect 5742 -4552 5798 -4496
rect 6132 -4544 6188 -4488
rect 6262 -4548 6318 -4492
rect 6652 -4542 6708 -4486
rect 6912 -4544 6968 -4488
rect 7042 -4542 7098 -4486
rect 7432 -4630 7488 -4574
rect 7562 -4628 7618 -4572
rect 8388 -4800 8484 -4704
rect 5036 -5056 5132 -4960
rect 12953 -3828 13207 -3574
rect 193 -5380 447 -5126
rect 5872 -5346 5928 -5290
rect 6002 -5348 6058 -5292
rect 6262 -5350 6318 -5294
rect 6652 -5348 6708 -5292
rect 6782 -5348 6838 -5292
rect 7172 -5352 7228 -5296
rect 7432 -5440 7488 -5384
rect 7562 -5438 7618 -5382
rect 8370 -5600 8466 -5504
rect 5032 -5856 5128 -5760
rect 193 -7080 447 -6826
rect 5032 -7044 5128 -6948
rect 5742 -6158 5798 -6102
rect 6002 -6146 6058 -6090
rect 6262 -6146 6318 -6090
rect 6652 -6142 6708 -6086
rect 6912 -6146 6968 -6090
rect 7172 -6138 7228 -6082
rect 7432 -6234 7488 -6178
rect 7562 -6238 7618 -6182
rect 6262 -6508 6318 -6452
rect 7300 -6510 7360 -6450
rect 6392 -6598 6448 -6542
rect 7430 -6600 7490 -6540
rect 6522 -6688 6578 -6632
rect 7560 -6690 7620 -6630
rect 6652 -6778 6708 -6722
rect 7690 -6780 7750 -6720
rect 6262 -7114 6318 -7058
rect 6636 -7108 6692 -7052
rect 7158 -7060 7214 -7004
rect 7692 -7256 7748 -7200
rect 8394 -6399 8490 -6303
rect 8372 -7582 8468 -7486
rect 12953 -5528 13207 -5274
rect 12953 -7228 13207 -6974
rect 193 -8928 447 -8674
rect 12953 -8928 13207 -8674
<< metal3 >>
rect 188 3254 452 3259
rect 12948 3254 13212 3259
rect 183 3000 193 3254
rect 447 3000 457 3254
rect 12943 3000 12953 3254
rect 13207 3000 13217 3254
rect 188 2995 452 3000
rect 12948 2995 13212 3000
rect 4980 1980 7340 2100
rect 188 1674 452 1679
rect 183 1420 193 1674
rect 447 1420 457 1674
rect 188 1415 452 1420
rect 5060 1085 5180 1980
rect 12948 1526 13212 1531
rect 12943 1272 12953 1526
rect 13207 1272 13217 1526
rect 12948 1267 13212 1272
rect 5032 1080 5180 1085
rect 5032 984 5042 1080
rect 5138 984 5180 1080
rect 5032 979 5180 984
rect 5060 860 5180 979
rect 5060 734 5180 740
rect 6163 604 6229 607
rect 5740 602 6229 604
rect 5740 546 6168 602
rect 6224 546 6229 602
rect 5740 544 6229 546
rect 2680 400 5000 520
rect 5120 400 5126 520
rect 188 -26 452 -21
rect 183 -280 193 -26
rect 447 -280 457 -26
rect 5740 -57 5800 544
rect 6163 541 6229 544
rect 7037 604 7103 609
rect 7037 548 7042 604
rect 7098 548 7103 604
rect 7037 543 7103 548
rect 5867 458 5933 463
rect 5867 402 5872 458
rect 5928 402 5933 458
rect 5867 397 5933 402
rect 5870 33 5930 397
rect 6000 123 6060 324
rect 6130 213 6190 324
rect 6127 208 6193 213
rect 6127 152 6132 208
rect 6188 152 6193 208
rect 6127 147 6193 152
rect 5997 118 6063 123
rect 5997 62 6002 118
rect 6058 62 6063 118
rect 5997 57 6063 62
rect 5867 28 5933 33
rect 5867 -28 5872 28
rect 5928 -28 5933 28
rect 5867 -33 5933 -28
rect 5737 -62 5803 -57
rect 5737 -118 5742 -62
rect 5798 -118 5803 -62
rect 5737 -123 5803 -118
rect 5052 -160 5168 -155
rect 5052 -256 5062 -160
rect 5158 -256 5168 -160
rect 5052 -261 5168 -256
rect 188 -285 452 -280
rect 5022 -960 5138 -955
rect 5022 -1056 5032 -960
rect 5128 -1056 5138 -960
rect 5022 -1061 5138 -1056
rect 2680 -1300 5020 -1180
rect 5140 -1300 5146 -1180
rect 5740 -1287 5800 -123
rect 5870 -485 5930 -33
rect 5867 -490 5933 -485
rect 5867 -546 5872 -490
rect 5928 -546 5933 -490
rect 5867 -551 5933 -546
rect 5737 -1292 5803 -1287
rect 5737 -1348 5742 -1292
rect 5798 -1348 5803 -1292
rect 5737 -1353 5803 -1348
rect 188 -1726 452 -1721
rect 183 -1980 193 -1726
rect 447 -1980 457 -1726
rect 5042 -1760 5158 -1755
rect 5042 -1856 5052 -1760
rect 5148 -1856 5158 -1760
rect 5042 -1861 5158 -1856
rect 188 -1985 452 -1980
rect 5036 -2559 5152 -2554
rect 5036 -2655 5046 -2559
rect 5142 -2655 5152 -2559
rect 5036 -2660 5152 -2655
rect 5740 -2879 5800 -1353
rect 5870 -2081 5930 -551
rect 5867 -2086 5933 -2081
rect 5867 -2142 5872 -2086
rect 5928 -2142 5933 -2086
rect 6000 -2087 6060 57
rect 6130 -479 6190 147
rect 6127 -484 6193 -479
rect 6127 -540 6132 -484
rect 6188 -540 6193 -484
rect 6127 -545 6193 -540
rect 6130 -1285 6190 -545
rect 6127 -1290 6193 -1285
rect 6127 -1346 6132 -1290
rect 6188 -1346 6193 -1290
rect 6127 -1351 6193 -1346
rect 5867 -2147 5933 -2142
rect 5997 -2092 6063 -2087
rect 2680 -3000 5020 -2880
rect 5140 -3000 5146 -2880
rect 5737 -2884 5803 -2879
rect 5737 -2940 5742 -2884
rect 5798 -2940 5803 -2884
rect 5737 -2945 5803 -2940
rect 5052 -3360 5168 -3355
rect 188 -3426 452 -3421
rect 183 -3680 193 -3426
rect 447 -3680 457 -3426
rect 5052 -3456 5062 -3360
rect 5158 -3456 5168 -3360
rect 5052 -3461 5168 -3456
rect 188 -3685 452 -3680
rect 5026 -4160 5142 -4155
rect 5026 -4256 5036 -4160
rect 5132 -4256 5142 -4160
rect 5026 -4261 5142 -4256
rect 5740 -4491 5800 -2945
rect 5870 -3679 5930 -2147
rect 5997 -2148 6002 -2092
rect 6058 -2148 6063 -2092
rect 5997 -2153 6063 -2148
rect 6000 -2881 6060 -2153
rect 5997 -2886 6063 -2881
rect 5997 -2942 6002 -2886
rect 6058 -2942 6063 -2886
rect 5997 -2947 6063 -2942
rect 5867 -3684 5933 -3679
rect 5867 -3740 5872 -3684
rect 5928 -3740 5933 -3684
rect 5867 -3745 5933 -3740
rect 5737 -4496 5803 -4491
rect 5737 -4552 5742 -4496
rect 5798 -4552 5803 -4496
rect 5737 -4557 5803 -4552
rect 2620 -4700 5020 -4580
rect 5140 -4700 5146 -4580
rect 5026 -4960 5142 -4955
rect 5026 -5056 5036 -4960
rect 5132 -5056 5142 -4960
rect 5026 -5061 5142 -5056
rect 188 -5126 452 -5121
rect 183 -5380 193 -5126
rect 447 -5380 457 -5126
rect 188 -5385 452 -5380
rect 5022 -5760 5138 -5755
rect 5022 -5856 5032 -5760
rect 5128 -5856 5138 -5760
rect 5022 -5861 5138 -5856
rect 5740 -6097 5800 -4557
rect 5870 -5285 5930 -3745
rect 5867 -5290 5933 -5285
rect 6000 -5287 6060 -2947
rect 6130 -3683 6190 -1351
rect 6260 -3679 6320 324
rect 6390 -479 6450 324
rect 6387 -484 6453 -479
rect 6387 -540 6392 -484
rect 6448 -540 6453 -484
rect 6387 -545 6453 -540
rect 6390 -1283 6450 -545
rect 6387 -1288 6453 -1283
rect 6387 -1344 6392 -1288
rect 6448 -1344 6453 -1288
rect 6387 -1349 6453 -1344
rect 6390 -2083 6450 -1349
rect 6387 -2088 6453 -2083
rect 6387 -2144 6392 -2088
rect 6448 -2144 6453 -2088
rect 6387 -2149 6453 -2144
rect 6390 -2885 6450 -2149
rect 6387 -2890 6453 -2885
rect 6387 -2946 6392 -2890
rect 6448 -2946 6453 -2890
rect 6387 -2951 6453 -2946
rect 6127 -3688 6193 -3683
rect 6127 -3744 6132 -3688
rect 6188 -3744 6193 -3688
rect 6127 -3749 6193 -3744
rect 6257 -3684 6323 -3679
rect 6257 -3740 6262 -3684
rect 6318 -3740 6323 -3684
rect 6257 -3745 6323 -3740
rect 6130 -4483 6190 -3749
rect 6127 -4488 6193 -4483
rect 6260 -4487 6320 -3745
rect 6127 -4544 6132 -4488
rect 6188 -4544 6193 -4488
rect 6127 -4549 6193 -4544
rect 6257 -4492 6323 -4487
rect 6257 -4548 6262 -4492
rect 6318 -4548 6323 -4492
rect 5867 -5346 5872 -5290
rect 5928 -5346 5933 -5290
rect 5867 -5351 5933 -5346
rect 5997 -5292 6063 -5287
rect 5997 -5348 6002 -5292
rect 6058 -5348 6063 -5292
rect 5737 -6102 5803 -6097
rect 5737 -6158 5742 -6102
rect 5798 -6158 5803 -6102
rect 5737 -6163 5803 -6158
rect 2680 -6400 5020 -6280
rect 5140 -6400 5146 -6280
rect 5740 -6460 5800 -6163
rect 5870 -6460 5930 -5351
rect 5997 -5353 6063 -5348
rect 6000 -6085 6060 -5353
rect 5997 -6090 6063 -6085
rect 5997 -6146 6002 -6090
rect 6058 -6146 6063 -6090
rect 5997 -6151 6063 -6146
rect 6000 -6460 6060 -6151
rect 6130 -6460 6190 -4549
rect 6257 -4553 6323 -4548
rect 6260 -5289 6320 -4553
rect 6257 -5294 6323 -5289
rect 6257 -5350 6262 -5294
rect 6318 -5350 6323 -5294
rect 6257 -5355 6323 -5350
rect 6260 -6085 6320 -5355
rect 6257 -6090 6323 -6085
rect 6257 -6146 6262 -6090
rect 6318 -6146 6323 -6090
rect 6257 -6151 6323 -6146
rect 6260 -6447 6320 -6151
rect 6257 -6452 6323 -6447
rect 6257 -6508 6262 -6452
rect 6318 -6508 6323 -6452
rect 6257 -6513 6323 -6508
rect 188 -6826 452 -6821
rect 183 -7080 193 -6826
rect 447 -7080 457 -6826
rect 5022 -6948 5138 -6943
rect 5022 -7044 5032 -6948
rect 5128 -7044 5138 -6948
rect 5022 -7049 5138 -7044
rect 6260 -7053 6320 -6513
rect 6390 -6537 6450 -2951
rect 6387 -6542 6453 -6537
rect 6387 -6598 6392 -6542
rect 6448 -6598 6453 -6542
rect 6387 -6603 6453 -6598
rect 6390 -7050 6450 -6603
rect 6520 -6627 6580 324
rect 6650 -481 6710 324
rect 6780 -55 6840 250
rect 6910 35 6970 250
rect 7040 125 7100 543
rect 8406 536 8522 541
rect 8406 440 8416 536
rect 8512 440 8522 536
rect 8406 435 8522 440
rect 7501 374 7567 377
rect 7170 372 7567 374
rect 7170 316 7506 372
rect 7562 316 7567 372
rect 7170 314 7567 316
rect 7170 215 7230 314
rect 7501 311 7567 314
rect 7165 210 7235 215
rect 7165 150 7170 210
rect 7230 150 7235 210
rect 7165 145 7235 150
rect 7035 120 7105 125
rect 7035 60 7040 120
rect 7100 60 7105 120
rect 7035 55 7105 60
rect 6905 30 6975 35
rect 6905 -30 6910 30
rect 6970 -30 6975 30
rect 6905 -35 6975 -30
rect 6775 -60 6845 -55
rect 6775 -120 6780 -60
rect 6840 -120 6845 -60
rect 6775 -125 6845 -120
rect 6780 -479 6840 -125
rect 6647 -486 6713 -481
rect 6647 -542 6652 -486
rect 6708 -542 6713 -486
rect 6647 -547 6713 -542
rect 6777 -484 6843 -479
rect 6777 -540 6782 -484
rect 6838 -540 6843 -484
rect 6777 -545 6843 -540
rect 6650 -1283 6710 -547
rect 6647 -1288 6713 -1283
rect 6647 -1344 6652 -1288
rect 6708 -1344 6713 -1288
rect 6647 -1349 6713 -1344
rect 6650 -2077 6710 -1349
rect 6647 -2082 6713 -2077
rect 6647 -2138 6652 -2082
rect 6708 -2138 6713 -2082
rect 6780 -2087 6840 -545
rect 6910 -1287 6970 -35
rect 7040 -491 7100 55
rect 7037 -496 7103 -491
rect 7037 -552 7042 -496
rect 7098 -552 7103 -496
rect 7037 -557 7103 -552
rect 7040 -1281 7100 -557
rect 7037 -1286 7103 -1281
rect 6907 -1292 6973 -1287
rect 6907 -1348 6912 -1292
rect 6968 -1348 6973 -1292
rect 7037 -1342 7042 -1286
rect 7098 -1342 7103 -1286
rect 7037 -1347 7103 -1342
rect 6907 -1353 6973 -1348
rect 6647 -2143 6713 -2138
rect 6777 -2092 6843 -2087
rect 6650 -2883 6710 -2143
rect 6777 -2148 6782 -2092
rect 6838 -2148 6843 -2092
rect 6777 -2153 6843 -2148
rect 6647 -2888 6713 -2883
rect 6647 -2944 6652 -2888
rect 6708 -2944 6713 -2888
rect 6647 -2949 6713 -2944
rect 6650 -3685 6710 -2949
rect 6647 -3690 6713 -3685
rect 6780 -3689 6840 -2153
rect 6910 -2887 6970 -1353
rect 6907 -2892 6973 -2887
rect 6907 -2948 6912 -2892
rect 6968 -2948 6973 -2892
rect 6907 -2953 6973 -2948
rect 6647 -3746 6652 -3690
rect 6708 -3746 6713 -3690
rect 6647 -3751 6713 -3746
rect 6777 -3694 6843 -3689
rect 6777 -3750 6782 -3694
rect 6838 -3750 6843 -3694
rect 6650 -4481 6710 -3751
rect 6777 -3755 6843 -3750
rect 6647 -4486 6713 -4481
rect 6647 -4542 6652 -4486
rect 6708 -4542 6713 -4486
rect 6647 -4547 6713 -4542
rect 6650 -5287 6710 -4547
rect 6780 -5287 6840 -3755
rect 6910 -4483 6970 -2953
rect 7040 -3693 7100 -1347
rect 7170 -2089 7230 145
rect 7300 -485 7360 -90
rect 7297 -490 7363 -485
rect 7297 -546 7302 -490
rect 7358 -546 7363 -490
rect 7297 -551 7363 -546
rect 7300 -1285 7360 -551
rect 7297 -1290 7363 -1285
rect 7297 -1346 7302 -1290
rect 7358 -1346 7363 -1290
rect 7297 -1351 7363 -1346
rect 7300 -2083 7360 -1351
rect 7297 -2088 7363 -2083
rect 7167 -2094 7233 -2089
rect 7167 -2150 7172 -2094
rect 7228 -2150 7233 -2094
rect 7297 -2144 7302 -2088
rect 7358 -2144 7363 -2088
rect 7297 -2149 7363 -2144
rect 7167 -2155 7233 -2150
rect 7170 -2893 7230 -2155
rect 7300 -2879 7360 -2149
rect 7297 -2884 7363 -2879
rect 7167 -2898 7233 -2893
rect 7167 -2954 7172 -2898
rect 7228 -2954 7233 -2898
rect 7297 -2940 7302 -2884
rect 7358 -2940 7363 -2884
rect 7297 -2945 7363 -2940
rect 7167 -2959 7233 -2954
rect 7037 -3698 7103 -3693
rect 7037 -3754 7042 -3698
rect 7098 -3754 7103 -3698
rect 7037 -3759 7103 -3754
rect 7040 -4481 7100 -3759
rect 6907 -4488 6973 -4483
rect 6907 -4544 6912 -4488
rect 6968 -4544 6973 -4488
rect 6907 -4549 6973 -4544
rect 7037 -4486 7103 -4481
rect 7037 -4542 7042 -4486
rect 7098 -4542 7103 -4486
rect 7037 -4547 7103 -4542
rect 6647 -5292 6713 -5287
rect 6647 -5348 6652 -5292
rect 6708 -5348 6713 -5292
rect 6647 -5353 6713 -5348
rect 6777 -5292 6843 -5287
rect 6777 -5348 6782 -5292
rect 6838 -5348 6843 -5292
rect 6777 -5353 6843 -5348
rect 6650 -6081 6710 -5353
rect 6647 -6086 6713 -6081
rect 6647 -6142 6652 -6086
rect 6708 -6142 6713 -6086
rect 6647 -6147 6713 -6142
rect 6517 -6632 6583 -6627
rect 6517 -6688 6522 -6632
rect 6578 -6688 6583 -6632
rect 6517 -6693 6583 -6688
rect 6520 -6830 6580 -6693
rect 6650 -6717 6710 -6147
rect 6647 -6722 6713 -6717
rect 6647 -6778 6652 -6722
rect 6708 -6778 6713 -6722
rect 6647 -6783 6713 -6778
rect 6650 -6830 6710 -6783
rect 6780 -6830 6840 -5353
rect 6910 -6085 6970 -4549
rect 6907 -6090 6973 -6085
rect 6907 -6146 6912 -6090
rect 6968 -6146 6973 -6090
rect 6907 -6151 6973 -6146
rect 6910 -6830 6970 -6151
rect 7040 -6830 7100 -4547
rect 7170 -5291 7230 -2959
rect 7167 -5296 7233 -5291
rect 7167 -5352 7172 -5296
rect 7228 -5352 7233 -5296
rect 7167 -5357 7233 -5352
rect 7170 -6077 7230 -5357
rect 7167 -6082 7233 -6077
rect 7167 -6138 7172 -6082
rect 7228 -6138 7233 -6082
rect 7167 -6143 7233 -6138
rect 7170 -6830 7230 -6143
rect 7300 -6445 7360 -2945
rect 7430 -3767 7490 -90
rect 7560 -561 7620 -90
rect 7557 -566 7623 -561
rect 7557 -622 7562 -566
rect 7618 -622 7623 -566
rect 7557 -627 7623 -622
rect 7560 -1379 7620 -627
rect 7557 -1384 7623 -1379
rect 7557 -1440 7562 -1384
rect 7618 -1440 7623 -1384
rect 7557 -1445 7623 -1440
rect 7560 -2163 7620 -1445
rect 7557 -2168 7623 -2163
rect 7557 -2224 7562 -2168
rect 7618 -2224 7623 -2168
rect 7557 -2229 7623 -2224
rect 7560 -2977 7620 -2229
rect 7557 -2982 7623 -2977
rect 7557 -3038 7562 -2982
rect 7618 -3038 7623 -2982
rect 7557 -3043 7623 -3038
rect 7427 -3772 7493 -3767
rect 7560 -3771 7620 -3043
rect 7427 -3828 7432 -3772
rect 7488 -3828 7493 -3772
rect 7427 -3833 7493 -3828
rect 7557 -3776 7623 -3771
rect 7557 -3832 7562 -3776
rect 7618 -3832 7623 -3776
rect 7430 -4569 7490 -3833
rect 7557 -3837 7623 -3832
rect 7560 -4567 7620 -3837
rect 7427 -4574 7493 -4569
rect 7427 -4630 7432 -4574
rect 7488 -4630 7493 -4574
rect 7427 -4635 7493 -4630
rect 7557 -4572 7623 -4567
rect 7557 -4628 7562 -4572
rect 7618 -4628 7623 -4572
rect 7557 -4633 7623 -4628
rect 7430 -5379 7490 -4635
rect 7560 -5377 7620 -4633
rect 7427 -5384 7493 -5379
rect 7427 -5440 7432 -5384
rect 7488 -5440 7493 -5384
rect 7427 -5445 7493 -5440
rect 7557 -5382 7623 -5377
rect 7557 -5438 7562 -5382
rect 7618 -5438 7623 -5382
rect 7557 -5443 7623 -5438
rect 7430 -6173 7490 -5445
rect 7427 -6178 7493 -6173
rect 7560 -6177 7620 -5443
rect 7427 -6234 7432 -6178
rect 7488 -6234 7493 -6178
rect 7427 -6239 7493 -6234
rect 7557 -6182 7623 -6177
rect 7557 -6238 7562 -6182
rect 7618 -6238 7623 -6182
rect 7295 -6450 7365 -6445
rect 7295 -6510 7300 -6450
rect 7360 -6510 7365 -6450
rect 7295 -6515 7365 -6510
rect 7300 -6830 7360 -6515
rect 7430 -6535 7490 -6239
rect 7557 -6243 7623 -6238
rect 7425 -6540 7495 -6535
rect 7425 -6600 7430 -6540
rect 7490 -6600 7495 -6540
rect 7425 -6605 7495 -6600
rect 7430 -6830 7490 -6605
rect 7560 -6625 7620 -6243
rect 7555 -6630 7625 -6625
rect 7555 -6690 7560 -6630
rect 7620 -6690 7625 -6630
rect 7555 -6695 7625 -6690
rect 7153 -7002 7219 -6999
rect 7560 -7002 7620 -6695
rect 7690 -6715 7750 -90
rect 12948 -174 13212 -169
rect 12943 -428 12953 -174
rect 13207 -428 13217 -174
rect 12948 -433 13212 -428
rect 8376 -704 8492 -699
rect 8376 -800 8386 -704
rect 8482 -800 8492 -704
rect 8376 -805 8492 -800
rect 8388 -1504 8504 -1499
rect 8388 -1600 8398 -1504
rect 8494 -1600 8504 -1504
rect 8388 -1605 8504 -1600
rect 12948 -1874 13212 -1869
rect 12943 -2128 12953 -1874
rect 13207 -2128 13217 -1874
rect 12948 -2133 13212 -2128
rect 8386 -2304 8502 -2299
rect 8386 -2400 8396 -2304
rect 8492 -2400 8502 -2304
rect 8386 -2405 8502 -2400
rect 8370 -3104 8486 -3099
rect 8370 -3200 8380 -3104
rect 8476 -3200 8486 -3104
rect 8370 -3205 8486 -3200
rect 12948 -3574 13212 -3569
rect 12943 -3828 12953 -3574
rect 13207 -3828 13217 -3574
rect 12948 -3833 13212 -3828
rect 8360 -3904 8476 -3899
rect 8360 -4000 8370 -3904
rect 8466 -4000 8476 -3904
rect 8360 -4005 8476 -4000
rect 8378 -4704 8494 -4699
rect 8378 -4800 8388 -4704
rect 8484 -4800 8494 -4704
rect 8378 -4805 8494 -4800
rect 12948 -5274 13212 -5269
rect 8360 -5504 8476 -5499
rect 8360 -5600 8370 -5504
rect 8466 -5600 8476 -5504
rect 12943 -5528 12953 -5274
rect 13207 -5528 13217 -5274
rect 12948 -5533 13212 -5528
rect 8360 -5605 8476 -5600
rect 8384 -6303 8500 -6298
rect 8384 -6399 8394 -6303
rect 8490 -6399 8500 -6303
rect 8384 -6404 8500 -6399
rect 7685 -6720 7755 -6715
rect 7685 -6780 7690 -6720
rect 7750 -6780 7755 -6720
rect 7685 -6785 7755 -6780
rect 7153 -7004 7620 -7002
rect 6631 -7050 6697 -7047
rect 6390 -7052 6697 -7050
rect 6257 -7058 6323 -7053
rect 188 -7085 452 -7080
rect 6257 -7114 6262 -7058
rect 6318 -7114 6323 -7058
rect 6390 -7108 6636 -7052
rect 6692 -7108 6697 -7052
rect 7153 -7060 7158 -7004
rect 7214 -7060 7620 -7004
rect 7153 -7062 7620 -7060
rect 7153 -7065 7219 -7062
rect 6390 -7110 6697 -7108
rect 6631 -7113 6697 -7110
rect 6257 -7119 6323 -7114
rect 7690 -7195 7750 -6785
rect 12948 -6974 13212 -6969
rect 7687 -7200 7753 -7195
rect 7687 -7256 7692 -7200
rect 7748 -7256 7753 -7200
rect 12943 -7228 12953 -6974
rect 13207 -7228 13217 -6974
rect 12948 -7233 13212 -7228
rect 7687 -7261 7753 -7256
rect 8362 -7486 8478 -7481
rect 8362 -7582 8372 -7486
rect 8468 -7582 8478 -7486
rect 8362 -7587 8478 -7582
rect 2680 -8100 5020 -7980
rect 5140 -8100 5190 -7980
rect 188 -8674 452 -8669
rect 183 -8928 193 -8674
rect 447 -8928 457 -8674
rect 188 -8933 452 -8928
rect 5070 -9828 5190 -8100
rect 12948 -8674 13212 -8669
rect 12943 -8928 12953 -8674
rect 13207 -8928 13217 -8674
rect 12948 -8933 13212 -8928
rect 5070 -9948 7380 -9828
<< via3 >>
rect 193 3000 447 3254
rect 12953 3000 13207 3254
rect 193 1420 447 1674
rect 12953 1272 13207 1526
rect 5042 984 5138 1080
rect 5060 740 5180 860
rect 5000 400 5120 520
rect 193 -280 447 -26
rect 5062 -256 5158 -160
rect 5032 -1056 5128 -960
rect 5020 -1300 5140 -1180
rect 193 -1980 447 -1726
rect 5052 -1856 5148 -1760
rect 5046 -2655 5142 -2559
rect 5020 -3000 5140 -2880
rect 193 -3680 447 -3426
rect 5062 -3456 5158 -3360
rect 5036 -4256 5132 -4160
rect 5020 -4700 5140 -4580
rect 5036 -5056 5132 -4960
rect 193 -5380 447 -5126
rect 5032 -5856 5128 -5760
rect 5020 -6400 5140 -6280
rect 193 -7080 447 -6826
rect 5032 -7044 5128 -6948
rect 8416 440 8512 536
rect 9490 252 9610 372
rect 12953 -428 13207 -174
rect 8386 -800 8482 -704
rect 9490 -1448 9610 -1328
rect 8398 -1600 8494 -1504
rect 12953 -2128 13207 -1874
rect 8396 -2400 8492 -2304
rect 8380 -3200 8476 -3104
rect 9490 -3148 9610 -3028
rect 12953 -3828 13207 -3574
rect 8370 -4000 8466 -3904
rect 8388 -4800 8484 -4704
rect 9500 -4848 9620 -4728
rect 8370 -5600 8466 -5504
rect 12953 -5528 13207 -5274
rect 8394 -6399 8490 -6303
rect 9490 -6548 9610 -6428
rect 12953 -7228 13207 -6974
rect 8372 -7582 8468 -7486
rect 5020 -8100 5140 -7980
rect 193 -8928 447 -8674
rect 9500 -8248 9620 -8128
rect 12953 -8928 13207 -8674
<< metal4 >>
rect 80 3254 548 3624
rect 80 3000 193 3254
rect 447 3000 548 3254
rect 80 1674 548 3000
rect 80 1420 193 1674
rect 447 1420 548 1674
rect 80 -26 548 1420
rect 12846 3254 13314 3634
rect 12846 3000 12953 3254
rect 13207 3000 13314 3254
rect 12846 1526 13314 3000
rect 12846 1272 12953 1526
rect 13207 1272 13314 1526
rect 80 -280 193 -26
rect 447 -280 548 -26
rect 80 -1726 548 -280
rect 80 -1980 193 -1726
rect 447 -1980 548 -1726
rect 80 -3426 548 -1980
rect 80 -3680 193 -3426
rect 447 -3680 548 -3426
rect 80 -5126 548 -3680
rect 80 -5380 193 -5126
rect 447 -5380 548 -5126
rect 80 -6826 548 -5380
rect 80 -7080 193 -6826
rect 447 -7080 548 -6826
rect 80 -8674 548 -7080
rect 4854 1080 5322 1266
rect 4854 984 5042 1080
rect 5138 984 5322 1080
rect 4854 860 5322 984
rect 4854 740 5060 860
rect 5180 740 5322 860
rect 4854 520 5322 740
rect 4854 400 5000 520
rect 5120 400 5322 520
rect 4854 -160 5322 400
rect 4854 -256 5062 -160
rect 5158 -256 5322 -160
rect 4854 -960 5322 -256
rect 4854 -1056 5032 -960
rect 5128 -1056 5322 -960
rect 4854 -1180 5322 -1056
rect 4854 -1300 5020 -1180
rect 5140 -1300 5322 -1180
rect 4854 -1760 5322 -1300
rect 4854 -1856 5052 -1760
rect 5148 -1856 5322 -1760
rect 4854 -2559 5322 -1856
rect 4854 -2655 5046 -2559
rect 5142 -2655 5322 -2559
rect 4854 -2880 5322 -2655
rect 4854 -3000 5020 -2880
rect 5140 -3000 5322 -2880
rect 4854 -3360 5322 -3000
rect 4854 -3456 5062 -3360
rect 5158 -3456 5322 -3360
rect 4854 -4160 5322 -3456
rect 4854 -4256 5036 -4160
rect 5132 -4256 5322 -4160
rect 4854 -4580 5322 -4256
rect 4854 -4700 5020 -4580
rect 5140 -4700 5322 -4580
rect 4854 -4960 5322 -4700
rect 4854 -5056 5036 -4960
rect 5132 -5056 5322 -4960
rect 4854 -5760 5322 -5056
rect 4854 -5856 5032 -5760
rect 5128 -5856 5322 -5760
rect 4854 -6280 5322 -5856
rect 4854 -6400 5020 -6280
rect 5140 -6400 5322 -6280
rect 4854 -6948 5322 -6400
rect 4854 -7044 5032 -6948
rect 5128 -7044 5322 -6948
rect 4854 -7746 5322 -7044
rect 8186 536 8654 738
rect 8186 440 8416 536
rect 8512 440 8654 536
rect 8186 -704 8654 440
rect 8186 -800 8386 -704
rect 8482 -800 8654 -704
rect 8186 -1504 8654 -800
rect 8186 -1600 8398 -1504
rect 8494 -1600 8654 -1504
rect 8186 -2304 8654 -1600
rect 8186 -2400 8396 -2304
rect 8492 -2400 8654 -2304
rect 8186 -3104 8654 -2400
rect 8186 -3200 8380 -3104
rect 8476 -3200 8654 -3104
rect 8186 -3904 8654 -3200
rect 8186 -4000 8370 -3904
rect 8466 -4000 8654 -3904
rect 8186 -4704 8654 -4000
rect 8186 -4800 8388 -4704
rect 8484 -4800 8654 -4704
rect 8186 -5504 8654 -4800
rect 8186 -5600 8370 -5504
rect 8466 -5600 8654 -5504
rect 8186 -6303 8654 -5600
rect 8186 -6399 8394 -6303
rect 8490 -6399 8654 -6303
rect 8186 -7486 8654 -6399
rect 8186 -7582 8372 -7486
rect 8468 -7582 8654 -7486
rect 8186 -7646 8654 -7582
rect 9266 372 9734 754
rect 9266 252 9490 372
rect 9610 252 9734 372
rect 9266 -1328 9734 252
rect 9266 -1448 9490 -1328
rect 9610 -1448 9734 -1328
rect 9266 -3028 9734 -1448
rect 9266 -3148 9490 -3028
rect 9610 -3148 9734 -3028
rect 9266 -4728 9734 -3148
rect 9266 -4848 9500 -4728
rect 9620 -4848 9734 -4728
rect 9266 -6428 9734 -4848
rect 9266 -6548 9490 -6428
rect 9610 -6548 9734 -6428
rect 9266 -7746 9734 -6548
rect 4854 -7980 9734 -7746
rect 4854 -8100 5020 -7980
rect 5140 -8100 9734 -7980
rect 4854 -8128 9734 -8100
rect 4854 -8248 9500 -8128
rect 9620 -8248 9734 -8128
rect 4854 -8254 9734 -8248
rect 12846 -174 13314 1272
rect 12846 -428 12953 -174
rect 13207 -428 13314 -174
rect 12846 -1874 13314 -428
rect 12846 -2128 12953 -1874
rect 13207 -2128 13314 -1874
rect 12846 -3574 13314 -2128
rect 12846 -3828 12953 -3574
rect 13207 -3828 13314 -3574
rect 12846 -5274 13314 -3828
rect 12846 -5528 12953 -5274
rect 13207 -5528 13314 -5274
rect 12846 -6974 13314 -5528
rect 12846 -7228 12953 -6974
rect 13207 -7228 13314 -6974
rect 80 -8928 193 -8674
rect 447 -8928 548 -8674
rect 80 -10046 548 -8928
rect 12846 -8674 13314 -7228
rect 12846 -8928 12953 -8674
rect 13207 -8928 13314 -8674
rect 12846 -10046 13314 -8928
rect 80 -10514 13314 -10046
use sized_switch  sized_switch_0
timestamp 1683929354
transform 1 0 -260 0 1 -7010
box 920 -1090 4438 448
use sized_switch  sized_switch_1
timestamp 1683929354
transform 1 0 -260 0 1 1490
box 920 -1090 4438 448
use sized_switch  sized_switch_2
timestamp 1683929354
transform 1 0 -260 0 1 -210
box 920 -1090 4438 448
use sized_switch  sized_switch_3
timestamp 1683929354
transform 1 0 -260 0 1 -1910
box 920 -1090 4438 448
use sized_switch  sized_switch_4
timestamp 1683929354
transform 1 0 -260 0 1 -3610
box 920 -1090 4438 448
use sized_switch  sized_switch_5
timestamp 1683929354
transform 1 0 -260 0 1 -5310
box 920 -1090 4438 448
use sized_switch  sized_switch_6
timestamp 1683929354
transform 1 0 8210 0 1 -5458
box 920 -1090 4438 448
use sized_switch  sized_switch_7
timestamp 1683929354
transform 1 0 8210 0 1 -7158
box 920 -1090 4438 448
use sized_switch  sized_switch_8
timestamp 1683929354
transform 1 0 8210 0 1 -3758
box 920 -1090 4438 448
use sized_switch  sized_switch_9
timestamp 1683929354
transform 1 0 8210 0 1 -2058
box 920 -1090 4438 448
use sized_switch  sized_switch_10
timestamp 1683929354
transform 1 0 8210 0 1 -358
box 920 -1090 4438 448
use sized_switch  sized_switch_11
timestamp 1683929354
transform 1 0 8210 0 1 1342
box 920 -1090 4438 448
use sized_switch  sized_switch_12
timestamp 1683929354
transform 1 0 2210 0 1 -8858
box 920 -1090 4438 448
use sized_switch  sized_switch_13
timestamp 1683929354
transform 1 0 6010 0 1 -8858
box 920 -1090 4438 448
use sized_switch  sized_switch_14
timestamp 1683929354
transform 1 0 2120 0 1 3070
box 920 -1090 4438 448
use sized_switch  sized_switch_15
timestamp 1683929354
transform 1 0 5920 0 1 3070
box 920 -1090 4438 448
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5438 0 1 -3152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1662439860
transform 1 0 5438 0 1 -6352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1662439860
transform 1 0 5438 0 1 -1552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1662439860
transform 1 0 5438 0 1 -2352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1662439860
transform 1 0 5438 0 1 -752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1662439860
transform 1 0 5438 0 1 -3952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1662439860
transform 1 0 5438 0 1 -4752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1662439860
transform 1 0 7782 0 1 -6352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1662439860
transform 1 0 7782 0 1 -5552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_9
timestamp 1662439860
transform 1 0 7782 0 1 -4752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_10
timestamp 1662439860
transform 1 0 7782 0 1 -3952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_11
timestamp 1662439860
transform 1 0 7782 0 1 -3152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_12
timestamp 1662439860
transform 1 0 7782 0 1 -2352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_13
timestamp 1662439860
transform 1 0 7782 0 1 -1552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_14
timestamp 1662439860
transform 1 0 7782 0 1 -752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_15
timestamp 1662439860
transform 1 0 5438 0 1 -5552
box -38 -48 314 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8134 0 1 -752
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_2
timestamp 1662439860
transform 1 0 5270 0 1 -2352
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_3
timestamp 1662439860
transform 1 0 8134 0 1 -1552
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_4
timestamp 1662439860
transform 1 0 5270 0 1 -752
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_5
timestamp 1662439860
transform 1 0 5270 0 1 -1552
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_6
timestamp 1662439860
transform 1 0 5713 0 1 -7533
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_7
timestamp 1662439860
transform 1 0 5270 0 1 -3152
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_8
timestamp 1662439860
transform 1 0 5270 0 1 -3952
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_9
timestamp 1662439860
transform 1 0 5270 0 1 -4752
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_10
timestamp 1662439860
transform 1 0 5270 0 1 -5552
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_11
timestamp 1662439860
transform 1 0 5270 0 1 -6352
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_12
timestamp 1662439860
transform 1 0 5690 0 1 488
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_13
timestamp 1662439860
transform 1 0 7689 0 1 -7533
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_14
timestamp 1662439860
transform 1 0 8134 0 1 -6352
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_15
timestamp 1662439860
transform 1 0 8134 0 1 -5552
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_16
timestamp 1662439860
transform 1 0 8134 0 1 -4752
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_17
timestamp 1662439860
transform 1 0 8134 0 1 -3952
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_18
timestamp 1662439860
transform 1 0 8134 0 1 -3152
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_19
timestamp 1662439860
transform 1 0 8134 0 1 -2352
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_20
timestamp 1662439860
transform 1 0 7666 0 1 488
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_2  x1
timestamp 1683919673
transform 1 0 5790 0 1 -752
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x2
timestamp 1683919673
transform 1 0 5790 0 1 -1552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x3
timestamp 1683919673
transform 1 0 5790 0 1 -2352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x4
timestamp 1683919673
transform 1 0 5790 0 1 -3152
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x5
timestamp 1683919673
transform 1 0 5790 0 1 -3952
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x6
timestamp 1683919673
transform 1 0 5790 0 1 -4752
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x7
timestamp 1683919673
transform 1 0 5790 0 1 -5552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x8
timestamp 1683919673
transform 1 0 5790 0 1 -6352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x9
timestamp 1683919673
transform 1 0 6786 0 1 -6352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x10
timestamp 1683919673
transform 1 0 6786 0 1 -5552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x11
timestamp 1683919673
transform 1 0 6786 0 1 -4752
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x12
timestamp 1683919673
transform 1 0 6786 0 1 -3952
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x13
timestamp 1683919673
transform 1 0 6786 0 1 -3152
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x14
timestamp 1683919673
transform 1 0 6786 0 1 -2352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x15
timestamp 1683919673
transform 1 0 6786 0 1 -1552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x16
timestamp 1683919673
transform 1 0 6786 0 1 -752
box -38 -48 958 592
use sky130_fd_sc_hd__inv_8  x17 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6785 0 1 -7533
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x18
timestamp 1662439860
transform 1 0 5881 0 1 -7533
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x19
timestamp 1662439860
transform 1 0 6762 0 1 488
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x20
timestamp 1662439860
transform 1 0 5858 0 1 488
box -38 -48 866 592
<< labels >>
rlabel metal4 6000 -10500 7500 -10100 1 OUT
port 4 n
rlabel metal4 5000 500 5200 700 1 VDD
port 19 n
rlabel metal4 8300 -7300 8500 -7100 1 GND
port 20 n
rlabel metal2 -300 2400 -200 2500 1 SIG0
port 21 n
rlabel metal2 -300 800 -200 900 1 SIG1
port 22 n
rlabel metal2 -300 -900 -200 -800 1 SIG2
port 23 n
rlabel metal2 -300 -2600 -200 -2500 1 SIG3
port 24 n
rlabel metal2 -300 -4300 -200 -4200 1 SIG4
port 25 n
rlabel metal2 -300 -6000 -200 -5900 1 SIG5
port 26 n
rlabel metal2 -300 -7700 -200 -7600 1 SIG6
port 27 n
rlabel metal2 -300 -9500 -200 -9400 1 SIG7
port 28 n
rlabel metal2 13600 -9500 13700 -9400 1 SIG8
port 29 n
rlabel metal2 13600 -7800 13700 -7700 1 SIG9
port 30 n
rlabel metal2 13600 -6100 13700 -6000 1 SIG10
port 31 n
rlabel metal2 13600 -4400 13700 -4300 1 SIG11
port 32 n
rlabel metal2 13600 -2700 13700 -2600 1 SIG12
port 33 n
rlabel metal2 13600 -1000 13700 -900 1 SIG13
port 34 n
rlabel metal2 13600 700 13700 800 1 SIG14
port 35 n
rlabel metal2 13600 2400 13700 2500 1 SIG15
port 36 n
rlabel metal3 5740 240 5800 300 1 SEL0
port 37 n
rlabel metal3 6000 240 6060 300 1 SEL1
port 38 n
rlabel metal3 6260 240 6320 300 1 SEL2
port 39 n
rlabel metal3 6520 240 6580 300 1 SEL3
port 40 n
<< end >>
