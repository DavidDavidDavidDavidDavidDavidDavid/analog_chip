* NGSPICE file created from wrapper_flattened.ext - technology: sky130A

.subckt wrapper_flattened gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12]
+ gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[17]
+ gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5] gpio_analog[6]
+ gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10] gpio_noesd[11]
+ gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16] gpio_noesd[17]
+ gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6]
+ gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10] io_analog[1]
+ io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4] io_analog[5]
+ io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd2 vccd1 vdda2 vdda1
X0 a_41723_677112# constant_gm_fingers_0.Vout a_43834_677960# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=4.3e+12p pd=3.172e+07u as=7.25e+12p ps=5.348e+07u w=5e+06u l=1e+06u
X1 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X2 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=3.235e+13p pd=2.2294e+08u as=1.3679e+14p ps=1.00302e+09u w=5e+06u l=500000u
R0 vssd2 constant_gm_fingers_0.VSS sky130_fd_pr__res_generic_m3 w=7.55e+07u l=1e+07u
X3 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X4 analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y analog_mux_0.sky130_fd_sc_hd__inv_2_4.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=2.51e+13p pd=1.7004e+08u as=2.624e+14p ps=1.70496e+09u w=5e+06u l=150000u
X6 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=7.39e+13p pd=5.3956e+08u as=2.9e+13p ps=2.116e+08u w=5e+06u l=500000u
X7 a_24084_271906# a_24084_271906# analog_mux_0.SIG6 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.25e+12p pd=5.348e+07u as=9.6e+12p ps=6.5e+07u w=2.5e+06u l=500000u
X8 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=2.075e+13p pd=1.383e+08u as=0p ps=0u w=5e+06u l=150000u
X9 a_287394_343809# gpio_analog[4] a_287588_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X10 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X11 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.17928e+14p pd=5.06904e+09u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=1e+06u
X12 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[11] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.304e+14p pd=8.5216e+08u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X13 analog_mux_0.x1.A gpio_analog[3] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X14 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.82653e+14p ps=9.7052e+09u w=5e+06u l=150000u
X15 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.54e+13p ps=3.1816e+08u w=5e+06u l=500000u
X16 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X17 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X18 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X19 analog_mux_0.x1.D gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X20 analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X21 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X22 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X23 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X24 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X25 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X26 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X27 analog_mux_0.x1.D gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X28 a_42819_684860# io_analog[9] a_43026_690893# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=2.32e+13p pd=1.6928e+08u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X29 analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y analog_mux_0.sky130_fd_sc_hd__inv_2_5.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X30 io_analog[8] io_analog[8] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=2.14535e+14p ps=1.68384e+09u w=5e+07u l=200000u
X31 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.595e+13p ps=1.1638e+08u w=5e+06u l=500000u
X32 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X33 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=1.595e+13p pd=1.1638e+08u as=0p ps=0u w=5e+06u l=500000u
X34 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X35 a_287588_343809# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_1.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X36 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=2.555e+13p pd=1.8022e+08u as=0p ps=0u w=5e+06u l=1e+06u
X37 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X38 io_analog[8] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X39 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=1.595e+13p pd=1.1638e+08u as=0p ps=0u w=5e+06u l=500000u
X40 a_537154_685355# a_534722_685355# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X41 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X42 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X43 io_analog[9] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X44 a_287394_349409# analog_mux_0.x1.B a_287588_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X45 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X46 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X47 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.83e+13p ps=1.2732e+08u w=5e+06u l=1e+06u
X48 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X49 constant_gm_fingers_0.VSS gpio_analog[6] analog_mux_0.x1.D constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X50 constant_gm_fingers_0.VSS gpio_analog[4] analog_mux_0.x1.B constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X51 a_287144_347009# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X52 a_534722_685355# a_537154_685355# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X53 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X54 analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y analog_mux_0.sky130_fd_sc_hd__inv_2_1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X55 gpio_analog[13] gpio_analog[13] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=3.18606e+14p ps=2.87548e+09u w=5e+07u l=200000u
X56 constant_gm_fingers_0.VSS analog_mux_0.SIG6 a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+13p ps=1.6928e+08u w=5e+06u l=1e+06u
X57 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X58 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+13p ps=5.2976e+08u w=5e+06u l=500000u
X59 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_287144_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X60 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X61 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X62 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X63 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X64 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X65 a_288390_347809# gpio_analog[4] a_288584_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X66 analog_mux_0.sky130_fd_sc_hd__inv_2_2.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X67 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X68 a_287588_349409# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_4.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X69 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X70 analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y analog_mux_0.sky130_fd_sc_hd__inv_2_7.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X71 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X72 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[14] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X73 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X74 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X75 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X76 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X77 analog_mux_0.SIG6 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X78 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X79 vdda2 gpio_analog[13] gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X80 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X81 analog_mux_0.sky130_fd_sc_hd__inv_2_0.A analog_mux_0.x1.A a_287588_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X82 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X83 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X84 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X85 vccd2 io_analog[9] io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X86 a_287588_347809# analog_mux_0.x1.B a_287394_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X87 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X88 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.74e+13p pd=1.2696e+08u as=0p ps=0u w=5e+06u l=1e+06u
X89 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X90 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X91 a_288584_347809# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X92 a_287394_345409# analog_mux_0.x1.C a_287144_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X93 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X94 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X95 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_0.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X96 gpio_analog[13] gpio_analog[13] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X97 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X98 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X99 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X100 analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X101 io_analog[0] io_analog[0] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=3.81686e+14p ps=3.65032e+09u w=5e+07u l=200000u
X102 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X103 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X104 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X105 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X106 analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y analog_mux_0.sky130_fd_sc_hd__inv_2_14.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X107 vdda1 a_536916_284434# analog_mux_0.SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X108 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X109 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X110 a_288390_343809# analog_mux_0.x1.C a_288140_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X111 analog_mux_0.x1.C gpio_analog[5] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X112 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X113 a_42819_684860# io_analog[8] a_40125_693523# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X114 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.685e+13p ps=3.2874e+08u w=5e+06u l=500000u
X115 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X116 vccd2 io_analog[8] io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X117 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_0.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 vccd1 io_analog[0] io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X119 io_analog[9] io_analog[9] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X120 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X121 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=1e+06u
R1 vssa2 constant_gm_fingers_0.VSS sky130_fd_pr__res_generic_m3 w=7.45e+07u l=2.6e+06u
X122 gpio_analog[12] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X123 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X124 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X125 vdda2 gpio_analog[5] analog_mux_0.x1.C vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X126 vdda2 gpio_analog[3] analog_mux_0.x1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X127 analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y analog_mux_0.sky130_fd_sc_hd__inv_2_11.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X128 a_287144_343809# gpio_analog[5] a_287394_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X129 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X130 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X131 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 constant_gm_fingers_0.VSS gpio_analog[5] analog_mux_0.x1.C constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X133 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X134 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_9.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X136 io_analog[0] io_analog[0] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X137 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X138 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X139 analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X140 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X141 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X142 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X143 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X144 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X145 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X146 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X147 a_288390_349409# gpio_analog[5] a_288140_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X148 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X149 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X150 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X151 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[7] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X152 analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X153 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X154 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X155 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X156 a_17579_272227# gpio_analog[12] analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.395e+13p ps=9.558e+07u w=5e+06u l=500000u
X157 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X158 io_analog[8] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X159 vccd1 io_analog[0] io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X160 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X161 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X162 analog_mux_0.x1.A gpio_analog[3] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X163 constant_gm_fingers_0.VSS gpio_analog[6] a_288140_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X164 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X165 a_530722_289355# analog_mux_0.SIG14 constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X166 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X167 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 gpio_analog[12] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X169 vdda2 a_24084_271906# analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X170 a_287144_349409# analog_mux_0.x1.C a_287394_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X171 gpio_analog[13] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X172 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[7] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X173 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_9.A analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X174 analog_mux_0.sky130_fd_sc_hd__inv_2_11.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X175 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X176 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X177 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X178 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X179 gpio_analog[12] gpio_analog[12] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X180 io_analog[0] io_analog[0] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X181 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X182 a_288140_347809# analog_mux_0.x1.C a_288390_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X183 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X184 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X185 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X187 a_288584_346209# analog_mux_0.x1.B a_288390_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X188 constant_gm_fingers_0.VSS gpio_analog[6] analog_mux_0.x1.D constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X189 constant_gm_fingers_0.VSS gpio_analog[4] analog_mux_0.x1.B constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X190 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X191 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[11] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X192 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[16] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X193 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X194 vdda2 gpio_analog[13] gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X195 a_288140_344609# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X196 a_540916_680434# a_540371_681998# a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X197 a_537154_685355# io_analog[1] a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.406e+07u as=0p ps=0u w=5e+06u l=500000u
X198 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_0.A analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X199 analog_mux_0.x1.B gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X200 analog_mux_0.SIG5 gpio_analog[12] a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X201 gpio_analog[13] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X202 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X203 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X204 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[11] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X207 a_536916_284434# analog_mux_0.SIG13 a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X208 analog_mux_0.x1.B gpio_analog[4] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X209 analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y analog_mux_0.sky130_fd_sc_hd__inv_2_3.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X210 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X211 vdda1 a_536916_284434# analog_mux_0.SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X213 gpio_analog[13] gpio_analog[13] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X214 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X215 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X216 vccd2 a_43834_677960# a_43834_677960# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X217 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+13p ps=4.232e+08u w=5e+06u l=500000u
X218 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X219 analog_mux_0.SIG7 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X220 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X221 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X222 analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[3] a_288584_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X223 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X225 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.83e+13p pd=1.2732e+08u as=0p ps=0u w=5e+06u l=150000u
X226 io_analog[1] io_analog[1] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X227 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X228 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X229 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X230 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[15] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X231 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X232 a_287144_348609# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X233 analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y analog_mux_0.sky130_fd_sc_hd__inv_2_6.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X234 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X235 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X236 vdda1 gpio_analog[1] gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.81686e+14p pd=3.65032e+09u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X237 analog_mux_0.SIG13 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.105e+13p pd=7.674e+07u as=0p ps=0u w=1.25e+06u l=1e+06u
X238 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X239 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X240 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X241 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X242 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X243 a_17579_272227# gpio_analog[12] analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X244 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X245 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG6 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X246 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X247 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X248 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X249 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X250 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X251 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X252 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X253 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_5.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X254 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X255 analog_mux_0.sky130_fd_sc_hd__inv_2_2.A analog_mux_0.x1.A a_287588_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X256 vccd1 io_analog[1] io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X257 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X258 a_41723_677112# constant_gm_fingers_0.Vout a_43834_677960# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X259 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X260 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X261 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X262 gpio_analog[1] gpio_analog[1] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X263 analog_mux_0.SIG7 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X264 a_287394_345409# gpio_analog[4] a_287588_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X265 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X266 vdda2 gpio_analog[12] gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X267 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_2.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X268 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X269 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X270 io_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X271 a_17579_272227# analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X272 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X273 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X274 analog_mux_0.sky130_fd_sc_hd__inv_2_5.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X275 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X276 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X277 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X278 gpio_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X279 constant_gm_fingers_0.VSS gpio_analog[6] a_287144_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X280 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X281 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X282 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X283 analog_mux_0.x1.A gpio_analog[3] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X284 a_288390_343809# analog_mux_0.x1.B a_288584_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X285 gpio_analog[12] gpio_analog[12] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X286 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X287 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X288 a_287588_345409# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_6.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X289 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_2.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X290 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X291 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X292 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X293 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y analog_mux_0.SIG14 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X294 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X295 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X296 analog_mux_0.SIG14 gpio_analog[1] a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X297 a_17579_272227# analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X298 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X299 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X300 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X301 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X302 analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y analog_mux_0.sky130_fd_sc_hd__inv_2_13.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X303 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X304 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X305 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X306 a_287588_343809# gpio_analog[4] a_287394_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X307 a_17579_272227# gpio_analog[12] analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X308 vdda2 gpio_analog[12] gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X309 constant_gm_fingers_0.VSS gpio_analog[3] analog_mux_0.x1.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X310 a_288584_343809# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X311 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X312 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X313 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_287144_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X314 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X315 vdda2 gpio_analog[6] analog_mux_0.x1.D vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X317 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X318 io_analog[10] constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.406e+07u as=0p ps=0u w=5e+06u l=1e+06u
X319 a_288390_349409# gpio_analog[4] a_288584_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X320 constant_gm_fingers_0.VSS gpio_analog[6] analog_mux_0.x1.D constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X321 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X322 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X323 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X324 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X325 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X326 a_540459_681940# io_analog[0] a_540271_687858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X327 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X328 analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X329 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X330 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X331 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout io_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X332 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X333 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[7] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X334 constant_gm_fingers_0.VSS a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X335 constant_gm_fingers_0.VSS gpio_analog[6] a_288140_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X336 a_43026_690893# io_analog[9] a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X337 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X338 io_analog[1] io_analog[1] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X339 analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X340 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X341 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X342 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X343 a_287588_349409# analog_mux_0.x1.B a_287394_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X344 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X345 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X346 a_288584_349409# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X347 a_287394_347009# gpio_analog[5] a_287144_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X348 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X349 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X350 constant_gm_fingers_0.VSS a_41723_677112# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X351 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X352 vdda1 gpio_analog[1] gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X353 a_540916_680434# a_540916_680434# a_540371_681998# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.348e+07u w=2.5e+06u l=500000u
X354 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X355 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X356 analog_mux_0.sky130_fd_sc_hd__inv_2_9.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X357 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X358 a_288584_347809# gpio_analog[4] a_288390_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X359 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_2.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X360 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X361 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_7.A analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 a_288390_345409# gpio_analog[5] a_288140_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X363 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X364 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X365 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X366 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X367 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X368 constant_gm_fingers_0.Vout a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=4.35e+12p pd=3.174e+07u as=0p ps=0u w=5e+06u l=1e+06u
X369 a_29040_272091# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X370 vccd2 a_43834_677960# constant_gm_fingers_0.Vout vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X371 vccd1 io_analog[1] io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X372 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X373 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X374 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X375 analog_mux_0.SIG6 a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X376 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_2.A analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X377 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X378 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X379 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X380 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y analog_mux_0.SIG13 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X381 gpio_analog[1] gpio_analog[1] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X382 a_287144_345409# analog_mux_0.x1.C a_287394_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X383 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X384 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X385 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X386 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X387 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X388 a_537154_685355# io_analog[1] a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X389 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X390 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X391 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X392 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X393 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X394 a_24084_271906# analog_mux_0.SIG6 a_29040_272091# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X395 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X396 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X397 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_5.A analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X398 a_540459_681940# io_analog[0] a_540271_687858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X399 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X400 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X401 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X402 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X403 a_288140_343809# analog_mux_0.x1.C a_288390_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X404 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X405 a_43834_677960# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X406 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X407 io_analog[0] io_analog[0] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X408 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X409 a_40125_693523# io_analog[8] a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X410 vdda1 a_536916_284434# analog_mux_0.SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X411 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X412 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X413 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X414 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X415 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[15] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X416 analog_mux_0.SIG5 gpio_analog[12] a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X417 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X418 a_40125_693523# io_analog[8] a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X419 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X420 analog_mux_0.x1.C gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X421 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X422 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_11.A analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X424 a_17579_272227# gpio_analog[13] a_14374_271026# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X425 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X426 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X427 analog_mux_0.x1.C gpio_analog[5] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X428 vccd1 io_analog[0] io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X429 a_536459_285940# gpio_analog[0] a_536271_291858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X430 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X431 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X432 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X433 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X434 analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y analog_mux_0.sky130_fd_sc_hd__inv_2_1.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X435 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X436 a_288140_349409# gpio_analog[5] a_288390_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X437 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X438 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X439 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X440 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X441 constant_gm_fingers_0.VSS a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X442 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X443 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X444 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X445 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X446 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X447 gpio_analog[13] gpio_analog[13] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X448 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X449 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X450 io_analog[0] io_analog[0] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X451 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X452 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X453 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X454 constant_gm_fingers_0.VSS a_41723_677112# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X455 constant_gm_fingers_0.VSS gpio_analog[5] analog_mux_0.x1.C constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X456 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X457 a_288140_346209# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X458 io_analog[1] io_analog[1] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X459 a_287144_344609# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X460 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X461 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X462 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X463 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X464 a_42819_684860# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X465 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_11.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X466 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X467 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X468 constant_gm_fingers_0.VSS analog_mux_0.SIG6 a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X469 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X470 analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y analog_mux_0.sky130_fd_sc_hd__inv_2_4.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X471 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X472 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X473 vdda2 gpio_analog[13] gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X474 io_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X475 vdda1 gpio_analog[0] gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X476 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X477 a_29040_272091# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X478 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X479 analog_mux_0.x1.D gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X480 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X481 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X482 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X483 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X484 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X485 analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[3] a_288584_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X486 analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X487 analog_mux_0.x1.D gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X488 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.x1.A a_287588_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X489 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X490 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X491 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X492 gpio_analog[13] gpio_analog[13] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X493 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X494 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X495 analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y analog_mux_0.sky130_fd_sc_hd__inv_2_0.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X496 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X497 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y analog_mux_0.SIG14 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X498 constant_gm_fingers_0.VSS analog_mux_0.SIG6 a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X499 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X500 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X501 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X502 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_15.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X503 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X504 analog_mux_0.sky130_fd_sc_hd__inv_2_8.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X505 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X506 analog_mux_0.SIG14 gpio_analog[1] a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X507 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X508 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X509 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X510 vdda2 gpio_analog[13] gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X511 a_536459_285940# gpio_analog[0] a_536271_291858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X512 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X513 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X514 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X515 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_3.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X516 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X517 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X518 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X519 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X521 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X522 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X523 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X524 constant_gm_fingers_0.VSS a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X525 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X526 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X527 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X528 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X529 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X530 a_287394_348609# analog_mux_0.x1.C a_287144_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X531 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X532 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X533 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X534 a_287394_347009# analog_mux_0.x1.B a_287588_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X535 vdda2 gpio_analog[3] analog_mux_0.x1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X536 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y analog_mux_0.SIG15 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X537 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X538 analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y analog_mux_0.sky130_fd_sc_hd__inv_2_8.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X539 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X540 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X541 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X542 a_14374_271026# gpio_analog[13] a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X543 vdda2 a_24084_271906# analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X544 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X545 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X546 analog_mux_0.sky130_fd_sc_hd__inv_2_3.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X547 constant_gm_fingers_0.Vout a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X548 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X549 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X550 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X551 constant_gm_fingers_0.VSS gpio_analog[6] a_287144_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X552 a_29040_272091# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X553 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X554 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X555 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X556 constant_gm_fingers_0.Vout a_43834_677960# a_43834_677960# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.4192e+12p pd=1.168e+07u as=0p ps=0u w=2.5e+06u l=500000u
X557 vccd1 io_analog[0] io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X558 a_288390_345409# analog_mux_0.x1.B a_288584_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X559 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X560 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X561 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y analog_mux_0.SIG15 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X562 analog_mux_0.sky130_fd_sc_hd__inv_2_5.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X563 a_42819_684860# io_analog[8] a_40125_693523# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X564 a_287588_347009# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_0.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X565 a_41723_677112# constant_gm_fingers_0.Vout a_43834_677960# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X566 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X567 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y analog_mux_0.SIG6 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X568 gpio_analog[13] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X569 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X570 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X571 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X572 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X573 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X574 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X575 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_288140_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X576 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X577 analog_mux_0.SIG14 gpio_analog[1] a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X578 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X579 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X580 a_287588_345409# gpio_analog[4] a_287394_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X581 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X582 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X583 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X584 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X585 analog_mux_0.sky130_fd_sc_hd__inv_2_8.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X586 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X587 a_288584_345409# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X588 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X589 a_42819_684860# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X590 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X591 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X592 gpio_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X593 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y analog_mux_0.SIG13 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X594 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X595 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X596 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X597 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X598 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X599 a_537154_685355# a_534722_685355# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X600 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X601 vdda2 gpio_analog[4] analog_mux_0.x1.B vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X602 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X603 io_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X604 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X605 constant_gm_fingers_0.VSS gpio_analog[5] analog_mux_0.x1.C constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X606 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X607 constant_gm_fingers_0.VSS gpio_analog[3] analog_mux_0.x1.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X608 analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y analog_mux_0.sky130_fd_sc_hd__inv_2_11.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X609 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X610 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X611 a_288584_343809# analog_mux_0.x1.B a_288390_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X612 io_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X613 analog_mux_0.SIG14 a_530722_289355# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X614 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X615 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X616 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X617 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X618 a_534722_685355# a_537154_685355# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X619 gpio_analog[13] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X620 constant_gm_fingers_0.VSS gpio_analog[6] a_288140_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X621 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X622 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X623 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X624 analog_mux_0.SIG7 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X625 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X626 gpio_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X627 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X628 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X629 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X630 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X631 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X632 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X633 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X634 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X635 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X636 a_43834_677960# constant_gm_fingers_0.Vout a_41723_677112# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X637 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X638 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X639 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X640 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X641 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X642 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X643 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X644 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X645 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X646 a_29040_272091# analog_mux_0.SIG6 a_24084_271906# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X647 analog_mux_0.sky130_fd_sc_hd__inv_2_11.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X648 a_288584_349409# gpio_analog[4] a_288390_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X649 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X650 a_29040_272091# analog_mux_0.SIG6 a_24084_271906# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X651 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X652 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X653 a_288390_347009# analog_mux_0.x1.C a_288140_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X654 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X655 a_540371_681998# a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X656 io_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X657 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X658 a_288140_347809# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X659 a_540916_680434# a_540371_681998# a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X660 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X661 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X662 a_42819_684860# io_analog[9] a_43026_690893# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X663 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X664 gpio_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X665 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X666 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X667 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X668 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X669 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X670 a_287144_347009# gpio_analog[5] a_287394_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X671 vccd2 io_analog[9] io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X672 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X673 a_42819_684860# io_analog[9] a_43026_690893# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X674 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X675 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X676 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X677 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X678 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X679 a_17579_272227# analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X680 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X681 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X682 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_9.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X683 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X684 analog_mux_0.SIG7 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X685 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[3] a_288584_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X686 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X687 analog_mux_0.x1.B gpio_analog[4] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X688 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_3.A analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X689 a_288140_345409# gpio_analog[5] a_288390_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X690 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X691 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X692 a_537154_685355# io_analog[1] a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X693 analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y analog_mux_0.sky130_fd_sc_hd__inv_2_2.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X694 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X695 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X696 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X697 analog_mux_0.SIG6 a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X698 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X699 io_analog[10] constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X700 a_540459_681940# io_analog[0] a_540271_687858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X701 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X702 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X703 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X704 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X705 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X706 a_14374_271026# gpio_analog[13] a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X707 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X708 analog_mux_0.SIG14 gpio_analog[1] a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X709 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X710 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X711 analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X712 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X713 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X714 analog_mux_0.x1.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X715 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X716 gpio_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X717 io_analog[10] constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X718 a_536459_285940# gpio_analog[0] a_536271_291858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X719 analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y analog_mux_0.sky130_fd_sc_hd__inv_2_6.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X720 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_4.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X721 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[16] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X722 io_analog[9] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X723 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X724 analog_mux_0.x1.D gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X726 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X727 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X728 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X729 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X730 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X731 a_287394_348609# analog_mux_0.x1.B a_287588_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X732 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X733 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X734 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X735 a_287144_346209# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X736 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X737 a_17579_272227# analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X738 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X739 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X740 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X741 analog_mux_0.sky130_fd_sc_hd__inv_2_4.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X742 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X743 a_42819_684860# io_analog[8] a_40125_693523# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X744 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y analog_mux_0.SIG6 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X745 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X746 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X747 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X748 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X749 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X750 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X751 analog_mux_0.SIG5 a_11871_265693# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X752 a_287588_348609# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_2.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X753 io_analog[8] io_analog[8] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X754 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X755 vccd2 io_analog[9] io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X756 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X757 a_17579_272227# gpio_analog[13] a_14374_271026# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X758 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X759 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X760 a_11871_265693# analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X761 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X762 analog_mux_0.sky130_fd_sc_hd__inv_2_3.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X763 analog_mux_0.sky130_fd_sc_hd__inv_2_5.A analog_mux_0.x1.A a_287588_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
R2 constant_gm_fingers_0.VSS vssd1 sky130_fd_pr__res_generic_m3 w=7.7e+07u l=5e+06u
X764 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X765 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y analog_mux_0.SIG6 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X766 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X768 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X769 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X770 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X771 a_287394_344609# gpio_analog[5] a_287144_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X772 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X773 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X774 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_5.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X775 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X776 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X777 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X778 analog_mux_0.sky130_fd_sc_hd__inv_2_10.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X779 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X780 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X781 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X782 vccd2 io_analog[8] io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X783 analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y analog_mux_0.sky130_fd_sc_hd__inv_2_13.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X784 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[14] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X785 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X786 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X787 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 a_43834_677960# constant_gm_fingers_0.Vout a_41723_677112# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X789 a_43026_690893# io_analog[9] a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X790 a_14374_271026# gpio_analog[13] a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X791 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X792 constant_gm_fingers_0.VSS gpio_analog[6] analog_mux_0.x1.D constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X793 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X794 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X795 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X796 vdda1 a_536916_284434# analog_mux_0.SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X797 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X798 analog_mux_0.SIG14 a_530722_289355# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X799 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X800 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X801 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X802 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X803 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X804 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X805 analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y analog_mux_0.sky130_fd_sc_hd__inv_2_10.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X806 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X807 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X808 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X809 analog_mux_0.SIG13 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X810 a_540459_681940# io_analog[0] a_540271_687858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X811 a_37693_693523# a_40125_693523# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X812 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_8.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X813 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X814 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X815 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 constant_gm_fingers_0.VSS gpio_analog[6] a_287144_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X817 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X818 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X819 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X820 vdda2 gpio_analog[5] analog_mux_0.x1.C vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X821 a_288390_348609# gpio_analog[5] a_288140_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X822 vdda1 a_536916_284434# analog_mux_0.SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X823 a_288390_347009# gpio_analog[4] a_288584_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X824 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X825 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X826 analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X827 io_analog[9] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X828 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X829 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X830 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X831 io_analog[9] io_analog[9] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X832 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X833 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X834 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X835 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X836 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X837 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_288140_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X838 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X839 constant_gm_fingers_0.VSS analog_mux_0.SIG6 a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X840 a_287144_348609# analog_mux_0.x1.C a_287394_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X841 constant_gm_fingers_0.VSS a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X842 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X843 a_287588_347009# analog_mux_0.x1.B a_287394_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X844 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X845 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X846 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_8.A analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X847 analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X848 a_288584_347009# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X849 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X850 a_42819_684860# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X851 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X852 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X853 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X854 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X855 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X856 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_4.A analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X857 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout io_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X858 gpio_analog[0] gpio_analog[0] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X859 analog_mux_0.SIG6 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X860 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X861 a_14374_271026# gpio_analog[13] a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X862 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X863 a_288584_345409# analog_mux_0.x1.B a_288390_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X864 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X865 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X866 io_analog[8] io_analog[8] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X867 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_5.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X868 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X869 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X870 vccd2 io_analog[9] io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X871 a_536916_284434# analog_mux_0.SIG13 a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X872 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X873 a_288140_343809# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X874 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X875 vdda1 gpio_analog[0] gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X876 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_5.A analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X877 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X878 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X879 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X880 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X881 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X882 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_8.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X883 a_540371_681998# a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X884 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X885 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X886 a_536916_284434# analog_mux_0.SIG13 a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X887 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X888 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X889 analog_mux_0.x1.B gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X890 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X891 io_analog[8] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X892 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X893 vccd2 io_analog[8] io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X894 gpio_analog[0] gpio_analog[0] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X895 analog_mux_0.x1.C gpio_analog[5] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X896 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X897 vccd2 a_43834_677960# constant_gm_fingers_0.Vout vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X898 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[16] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X899 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_11.A analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X900 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[3] a_288584_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X901 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X902 a_43834_677960# constant_gm_fingers_0.Vout a_41723_677112# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X903 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X904 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X905 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X906 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X907 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X908 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X909 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X910 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X911 a_288140_349409# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X912 a_287144_347809# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X913 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X914 analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y analog_mux_0.sky130_fd_sc_hd__inv_2_15.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X915 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X916 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X917 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X918 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X919 vdda1 gpio_analog[0] gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X920 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[11] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X921 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X922 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X923 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X924 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X925 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X926 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X927 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X928 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X929 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X930 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X931 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X932 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X933 analog_mux_0.SIG5 a_11871_265693# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X934 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_11.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X935 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X936 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X937 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[3] a_288584_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X938 analog_mux_0.sky130_fd_sc_hd__inv_2_4.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X939 analog_mux_0.sky130_fd_sc_hd__inv_2_3.A analog_mux_0.x1.A a_287588_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X940 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X941 vccd2 a_43834_677960# a_43834_677960# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X942 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X943 gpio_analog[0] gpio_analog[0] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X944 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X945 a_288140_347009# analog_mux_0.x1.C a_288390_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X946 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X947 a_11871_265693# analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X948 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[15] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X949 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X950 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X951 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X952 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X953 vccd2 io_analog[8] io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X954 analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X955 a_540916_680434# a_540371_681998# a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X956 io_analog[9] io_analog[9] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X957 analog_mux_0.x1.D gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X958 a_287394_344609# gpio_analog[4] a_287588_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X959 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X960 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X961 a_536916_284434# analog_mux_0.SIG13 a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X962 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X963 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X964 a_42819_684860# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X965 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X966 analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X967 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X968 a_43026_690893# io_analog[9] a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X969 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X970 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X971 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X972 analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y analog_mux_0.sky130_fd_sc_hd__inv_2_0.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X973 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X974 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X975 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X976 a_17579_272227# gpio_analog[13] a_14374_271026# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X977 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X978 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X979 a_287588_344609# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_15.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X980 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X981 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X982 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[14] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X983 a_42819_684860# io_analog[8] a_40125_693523# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X984 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X985 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X986 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X987 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X988 io_analog[8] io_analog[8] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X989 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X990 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X991 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X992 io_analog[8] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X993 gpio_analog[1] gpio_analog[1] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X994 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X995 a_37693_693523# a_40125_693523# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X996 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X997 vdda2 a_24084_271906# analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X998 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X999 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1000 constant_gm_fingers_0.VSS gpio_analog[6] a_287144_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1001 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1002 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1003 io_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1004 vdda2 gpio_analog[3] analog_mux_0.x1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1005 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1006 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1007 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1008 a_288390_348609# gpio_analog[4] a_288584_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X1009 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1010 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1011 a_42819_684860# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1012 analog_mux_0.sky130_fd_sc_hd__inv_2_4.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1013 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1014 constant_gm_fingers_0.VSS gpio_analog[3] analog_mux_0.x1.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1015 analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y analog_mux_0.sky130_fd_sc_hd__inv_2_8.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1016 gpio_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1017 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1018 gpio_analog[12] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1019 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y analog_mux_0.SIG14 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1020 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1021 vdda1 gpio_analog[1] gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1022 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1023 analog_mux_0.sky130_fd_sc_hd__inv_2_5.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1024 a_287588_348609# analog_mux_0.x1.B a_287394_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1025 a_288584_348609# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1026 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1027 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1028 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1029 a_287394_346209# analog_mux_0.x1.C a_287144_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X1030 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1031 analog_mux_0.x1.B gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1032 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_3.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1034 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1035 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1036 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1037 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1038 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1039 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1040 io_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1041 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1042 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1043 analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1045 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1046 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout io_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1047 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1048 a_288390_344609# analog_mux_0.x1.C a_288140_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X1049 analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1050 gpio_analog[0] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1051 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y gpio_analog[7] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1052 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1053 vdda2 gpio_analog[4] analog_mux_0.x1.B vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1055 analog_mux_0.SIG7 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1056 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1057 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_3.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1058 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout io_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1059 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1060 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R3 constant_gm_fingers_0.VSS vssa1 sky130_fd_pr__res_generic_m4 w=2.75e+07u l=2.8e+06u
X1061 constant_gm_fingers_0.VSS gpio_analog[4] analog_mux_0.x1.B constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1062 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1063 a_17579_272227# analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1064 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_3.A analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1065 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1066 analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y analog_mux_0.sky130_fd_sc_hd__inv_2_12.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1067 a_287144_344609# gpio_analog[5] a_287394_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1068 a_540916_680434# a_540371_681998# a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1069 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1070 a_537154_685355# io_analog[1] a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1071 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1072 io_analog[8] io_analog[8] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1073 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_10.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1074 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1075 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1076 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1077 a_536916_284434# analog_mux_0.SIG13 a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1078 a_540459_681940# io_analog[0] a_540271_687858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1079 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG6 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1080 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1081 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1082 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1083 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1084 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1085 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1086 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1087 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1088 vdda2 gpio_analog[12] gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1089 vccd1 io_analog[1] io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1090 constant_gm_fingers_0.Vout a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1091 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1092 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_288140_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1093 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1094 gpio_analog[1] gpio_analog[1] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1095 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1096 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1097 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_10.A analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1100 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1101 a_17579_272227# analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1102 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1103 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_13.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1104 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1105 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1106 vccd1 io_analog[1] io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1107 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1108 analog_mux_0.x1.C gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1109 a_288140_348609# gpio_analog[5] a_288390_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1110 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1111 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1112 a_288584_347009# gpio_analog[4] a_288390_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1113 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1114 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1115 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1116 io_analog[1] io_analog[1] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1117 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1118 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1119 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1120 a_40125_693523# a_37693_693523# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X1121 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1122 analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1123 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1124 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1125 analog_mux_0.SIG6 a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1126 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y gpio_analog[15] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1127 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1128 a_288140_345409# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1129 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1130 a_287144_343809# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1131 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1132 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1133 vdda1 gpio_analog[1] gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1134 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1135 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1136 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1137 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1138 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1139 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 a_537154_685355# io_analog[1] a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1141 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1142 analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y analog_mux_0.sky130_fd_sc_hd__inv_2_2.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1143 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1144 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1145 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1146 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1147 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1148 analog_mux_0.x1.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1149 analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[3] a_288584_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1150 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1151 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1152 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1153 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.x1.A a_287588_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1154 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1155 analog_mux_0.x1.A gpio_analog[3] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1156 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1157 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1158 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1159 a_287144_349409# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1160 analog_mux_0.x1.D gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1161 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1162 analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y analog_mux_0.sky130_fd_sc_hd__inv_2_5.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1163 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1164 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1165 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1166 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1167 analog_mux_0.SIG14 gpio_analog[1] a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1168 gpio_analog[0] gpio_analog[0] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1169 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1170 analog_mux_0.x1.D gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1171 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1172 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1173 a_536459_285940# gpio_analog[0] a_536271_291858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1174 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1175 vdda2 gpio_analog[6] analog_mux_0.x1.D vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1176 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1177 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1178 vdda2 gpio_analog[4] analog_mux_0.x1.B vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1179 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1180 vdda1 gpio_analog[0] gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1181 analog_mux_0.sky130_fd_sc_hd__inv_2_4.A analog_mux_0.x1.A a_287588_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1182 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1183 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1184 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1185 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1186 a_43026_690893# io_analog[9] a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1187 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1188 a_43834_677960# a_43834_677960# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1189 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1190 vccd1 io_analog[1] io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1191 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1192 a_287394_347809# gpio_analog[5] a_287144_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1193 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y analog_mux_0.SIG14 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1194 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1195 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1196 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1197 a_287394_346209# gpio_analog[4] a_287588_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1198 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_4.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1199 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1200 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1201 gpio_analog[0] gpio_analog[0] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1202 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1203 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1204 analog_mux_0.sky130_fd_sc_hd__inv_2_0.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1205 gpio_analog[1] gpio_analog[1] vdda1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1206 io_analog[10] constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1207 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1208 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1209 vdda1 gpio_analog[1] gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1210 constant_gm_fingers_0.Vout constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X1211 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_287144_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1212 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1213 a_540916_680434# a_540916_680434# a_540371_681998# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1214 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1215 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1216 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1217 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1218 a_288390_344609# analog_mux_0.x1.B a_288584_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1219 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1220 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1221 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1222 analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1223 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 a_536916_284434# a_536916_284434# analog_mux_0.SIG13 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1225 a_287588_346209# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_5.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1226 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_4.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1227 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1228 a_24084_271906# analog_mux_0.SIG6 a_29040_272091# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1229 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1230 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1231 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1232 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1233 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1234 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1235 io_analog[1] io_analog[1] vccd1 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1236 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1237 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1238 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1239 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1240 analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y analog_mux_0.sky130_fd_sc_hd__inv_2_14.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1241 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1242 constant_gm_fingers_0.VSS analog_mux_0.SIG6 a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1243 a_287588_344609# gpio_analog[4] a_287394_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1244 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1245 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1246 analog_mux_0.SIG14 gpio_analog[1] a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1247 analog_mux_0.x1.C gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1248 a_288584_344609# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1249 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1250 io_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1251 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1253 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1254 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1255 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y analog_mux_0.SIG15 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1256 analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y analog_mux_0.sky130_fd_sc_hd__inv_2_10.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1257 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1258 a_24084_271906# analog_mux_0.SIG6 a_29040_272091# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1259 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1260 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1261 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1262 a_540459_681940# io_analog[0] a_540271_687858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1263 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1264 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1265 vdda2 gpio_analog[5] analog_mux_0.x1.C vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1266 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1267 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1268 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_288140_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1269 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1270 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1272 constant_gm_fingers_0.VSS analog_mux_0.SIG6 a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1273 analog_mux_0.sky130_fd_sc_hd__inv_2_3.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1274 constant_gm_fingers_0.VSS gpio_analog[5] analog_mux_0.x1.C constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1275 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1276 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1277 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1278 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1279 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1280 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1281 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y analog_mux_0.SIG13 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1282 analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1283 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1284 analog_mux_0.x1.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1285 analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 a_288584_348609# gpio_analog[4] a_288390_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1287 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1288 a_40125_693523# a_37693_693523# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X1289 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1290 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1291 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_4.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1292 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1293 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1294 a_43834_677960# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1295 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1296 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_8.A analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1297 a_288390_346209# gpio_analog[5] a_288140_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1298 vccd2 a_43834_677960# a_43834_677960# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1299 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1300 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1301 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1302 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1303 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1304 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1305 vdda1 gpio_analog[0] gpio_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1306 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1307 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1308 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1309 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_4.A analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1310 a_536916_284434# a_536916_284434# analog_mux_0.SIG13 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1311 vccd1 io_analog[0] io_analog[0] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1312 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1313 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1314 a_287144_346209# analog_mux_0.x1.C a_287394_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1315 vdda2 gpio_analog[6] analog_mux_0.x1.D vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1316 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1317 vdda2 gpio_analog[4] analog_mux_0.x1.B vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1318 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1319 a_540371_681998# a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1320 gpio_analog[12] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1321 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1322 constant_gm_fingers_0.VSS analog_mux_0.SIG6 a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1323 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A analog_mux_0.x1.C vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1324 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1326 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1327 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1328 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1329 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1330 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1331 analog_mux_0.SIG13 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1332 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1333 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1334 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1335 gpio_analog[8] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1336 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1337 analog_mux_0.SIG6 a_24084_271906# a_24084_271906# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1338 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_0.A analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1339 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1340 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1341 a_288140_344609# analog_mux_0.x1.C a_288390_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1342 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1343 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y gpio_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1344 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1345 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1346 analog_mux_0.x1.B gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1347 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1348 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1349 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1350 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1351 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1352 analog_mux_0.x1.B gpio_analog[4] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1353 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1354 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1355 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1356 gpio_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1357 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1358 vdda2 gpio_analog[13] gpio_analog[13] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1359 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1360 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1361 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1362 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1363 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1364 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1365 analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1366 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1367 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1368 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1369 io_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1370 gpio_analog[13] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1371 analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y analog_mux_0.sky130_fd_sc_hd__inv_2_15.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1372 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1373 a_42819_684860# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1374 constant_gm_fingers_0.VSS a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1375 a_536459_285940# gpio_analog[0] a_536271_291858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1376 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1377 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1378 analog_mux_0.SIG7 analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1379 gpio_analog[7] analog_mux_0.sky130_fd_sc_hd__inv_2_4.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1380 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1381 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1382 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1383 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1384 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1385 a_287394_347809# analog_mux_0.x1.B a_287588_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1386 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1387 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1388 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1389 a_288140_347009# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1390 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1391 a_287144_345409# gpio_analog[6] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1392 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1393 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1394 io_analog[9] io_analog[9] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1395 analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1396 analog_mux_0.sky130_fd_sc_hd__inv_2_2.A analog_mux_0.x1.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1397 a_29040_272091# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X1398 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1399 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1400 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1401 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_12.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1402 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1403 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1404 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1405 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1406 a_40125_693523# io_analog[8] a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1407 analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1408 a_29040_272091# analog_mux_0.SIG6 a_24084_271906# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1409 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1410 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1411 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1412 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1413 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1414 a_287588_347809# analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_3.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1415 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1416 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1417 io_analog[10] constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1418 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1419 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1420 io_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1421 analog_mux_0.sky130_fd_sc_hd__inv_2_11.A gpio_analog[3] a_288584_347009# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1422 analog_mux_0.sky130_fd_sc_hd__inv_2_0.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1423 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.x1.A a_287588_345409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1424 a_537154_685355# io_analog[1] a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1425 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1426 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_2.A gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1427 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1428 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1429 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1430 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1431 analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y analog_mux_0.sky130_fd_sc_hd__inv_2_3.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1432 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1433 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1434 analog_mux_0.x1.A gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1435 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1436 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1437 a_287394_343809# gpio_analog[5] a_287144_343809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1438 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1439 analog_mux_0.SIG14 gpio_analog[1] a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1440 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1441 analog_mux_0.SIG15 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1442 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y analog_mux_0.SIG15 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1443 vdda2 analog_mux_0.x1.A analog_mux_0.sky130_fd_sc_hd__inv_2_6.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1444 constant_gm_fingers_0.VSS a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1445 analog_mux_0.sky130_fd_sc_hd__inv_2_9.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1446 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1447 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1448 a_536459_285940# gpio_analog[0] a_536271_291858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1449 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1450 constant_gm_fingers_0.VSS a_41723_677112# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1451 analog_mux_0.SIG13 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1452 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.SIG15 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1453 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1454 a_540371_681998# a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1455 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1456 analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y analog_mux_0.sky130_fd_sc_hd__inv_2_12.A constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1457 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1458 gpio_analog[12] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1459 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1460 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1461 vdda2 gpio_analog[3] analog_mux_0.x1.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1463 analog_mux_0.sky130_fd_sc_hd__inv_2_4.A analog_mux_0.x1.D vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y analog_mux_0.SIG6 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1465 constant_gm_fingers_0.VSS gpio_analog[3] analog_mux_0.x1.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1466 gpio_analog[12] gpio_analog[12] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1467 analog_mux_0.SIG7 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1468 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_13.A analog_mux_0.SIG14 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1469 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1470 a_287394_349409# analog_mux_0.x1.C a_287144_349409# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1471 gpio_analog[15] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1472 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1473 vdda2 gpio_analog[6] analog_mux_0.x1.D vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1474 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1475 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1476 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1477 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1478 a_42819_684860# constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1479 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1480 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1481 analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y analog_mux_0.sky130_fd_sc_hd__inv_2_9.A vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1482 a_43834_677960# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1483 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1484 gpio_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1485 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1486 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1487 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1488 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y analog_mux_0.SIG13 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1489 vdda2 gpio_analog[12] gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1490 io_analog[9] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1491 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[14] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1492 constant_gm_fingers_0.VSS analog_mux_0.x1.D a_287144_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1493 constant_gm_fingers_0.Vout constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X1494 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1495 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1496 a_288390_347809# analog_mux_0.x1.C a_288140_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1497 a_288390_346209# analog_mux_0.x1.B a_288584_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1498 analog_mux_0.x1.B gpio_analog[4] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1499 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1500 analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1501 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1502 analog_mux_0.SIG5 gpio_analog[12] a_17579_272227# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1503 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1504 gpio_analog[12] gpio_analog[12] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1505 constant_gm_fingers_0.VSS gpio_analog[6] a_288140_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1506 gpio_analog[9] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1507 vdda1 a_536916_284434# analog_mux_0.SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1508 a_540916_680434# a_540371_681998# a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1509 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_15.A analog_mux_0.SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1510 a_287144_347809# gpio_analog[5] a_287394_347809# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1511 analog_mux_0.sky130_fd_sc_hd__inv_2_1.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1512 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1513 a_287588_346209# gpio_analog[4] a_287394_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1514 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1515 analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1516 gpio_analog[10] analog_mux_0.sky130_fd_sc_hd__inv_2_0.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1517 vdda2 gpio_analog[4] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 a_288584_346209# gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1519 constant_gm_fingers_0.VSS gpio_analog[4] analog_mux_0.x1.B constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1520 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1521 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1522 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_9.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1523 gpio_analog[16] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1524 vdda2 gpio_analog[12] gpio_analog[12] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1525 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1526 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_2.A analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 gpio_analog[1] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1528 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1529 a_540916_680434# a_540371_681998# a_541059_678436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1530 a_288584_344609# analog_mux_0.x1.B a_288390_344609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1531 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1532 vdda2 analog_mux_0.x1.C analog_mux_0.sky130_fd_sc_hd__inv_2_6.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1533 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1534 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1535 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1536 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1537 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1538 vdda2 gpio_analog[3] analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1539 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1540 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1541 a_537154_685355# io_analog[1] a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1542 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1543 gpio_analog[12] gpio_analog[12] vdda2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1544 analog_mux_0.SIG6 analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1545 io_analog[2] a_540371_681998# constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1546 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1547 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1548 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1549 analog_mux_0.SIG14 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1550 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1551 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1552 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_12.A analog_mux_0.SIG13 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1553 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1554 constant_gm_fingers_0.VSS a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X1555 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_6.A analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1556 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1557 constant_gm_fingers_0.VSS a_41723_677112# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1558 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_8.A gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1559 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1560 a_540459_681940# io_analog[0] a_540271_687858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1561 vdda1 a_536271_291858# analog_mux_0.SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1562 a_17579_272227# analog_mux_0.SIG6 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1563 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1564 io_analog[8] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1565 constant_gm_fingers_0.VSS analog_mux_0.SIG13 a_536459_285940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1566 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout a_42819_684860# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1567 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1568 vdda2 analog_mux_0.x1.B analog_mux_0.sky130_fd_sc_hd__inv_2_7.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS gpio_analog[1] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1570 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1571 analog_mux_0.sky130_fd_sc_hd__inv_2_12.A gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1572 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_1.A analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1573 a_536459_285940# gpio_analog[0] a_536271_291858# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1574 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1575 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout io_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1576 a_530722_289355# analog_mux_0.SIG14 constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X1577 constant_gm_fingers_0.VSS analog_mux_0.sky130_fd_sc_hd__inv_2_10.A analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1578 constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1579 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1580 vdda2 a_14374_271026# analog_mux_0.SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1581 vdda2 analog_mux_0.SIG5 analog_mux_0.SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1582 analog_mux_0.x1.C gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1583 a_288140_348609# analog_mux_0.x1.D constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1584 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1585 analog_mux_0.SIG5 analog_mux_0.sky130_fd_sc_hd__inv_2_6.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1586 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y gpio_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1587 analog_mux_0.x1.C gpio_analog[5] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1588 constant_gm_fingers_0.VSS constant_gm_fingers_0.Vout io_analog[10] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1589 analog_mux_0.SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1590 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1591 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_3.A gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1592 gpio_analog[11] analog_mux_0.sky130_fd_sc_hd__inv_2_5.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1593 vdda2 gpio_analog[5] analog_mux_0.sky130_fd_sc_hd__inv_2_14.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1594 analog_mux_0.SIG7 analog_mux_0.SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1595 vdda1 analog_mux_0.SIG14 analog_mux_0.SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1596 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1597 vdda2 analog_mux_0.sky130_fd_sc_hd__inv_2_7.A analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1598 io_analog[10] constant_gm_fingers_0.Vout constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1599 constant_gm_fingers_0.VSS a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X1600 analog_mux_0.SIG15 analog_mux_0.sky130_fd_sc_hd__inv_2_14.A gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1601 gpio_analog[14] analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y gpio_analog[2] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1602 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1603 vdda2 gpio_analog[5] analog_mux_0.x1.C vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 vccd2 io_analog[9] io_analog[9] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1605 io_analog[9] constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1606 vdda2 gpio_analog[6] analog_mux_0.sky130_fd_sc_hd__inv_2_10.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1607 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_9.A constant_gm_fingers_0.VSS vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1608 vdda2 analog_mux_0.x1.D analog_mux_0.sky130_fd_sc_hd__inv_2_15.A vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 analog_mux_0.SIG13 analog_mux_0.SIG13 constant_gm_fingers_0.VSS constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1610 gpio_analog[2] analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y gpio_analog[16] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1611 analog_mux_0.sky130_fd_sc_hd__inv_2_13.A gpio_analog[3] a_288584_348609# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1612 analog_mux_0.sky130_fd_sc_hd__inv_2_2.A analog_mux_0.x1.B vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1613 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1614 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1615 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1616 vccd2 io_analog[8] io_analog[8] constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1617 constant_gm_fingers_0.VSS analog_mux_0.SIG6 analog_mux_0.SIG7 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1618 a_17579_272227# gpio_analog[12] analog_mux_0.SIG5 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1619 a_288140_346209# gpio_analog[5] a_288390_346209# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1620 io_analog[9] io_analog[9] vccd2 constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1621 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1622 a_536916_284434# analog_mux_0.SIG13 a_537059_282436# constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1623 vccd2 a_43834_677960# constant_gm_fingers_0.Vout vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

