* NGSPICE file created from lvs.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_UXPKRJ a_n621_n5174# a_114_n5088# a_n29_n5000# a_n474_n5088#
+ a_n323_n5000# a_461_n5000# a_167_n5000# a_69_n5000# a_16_5022# a_310_n5088# a_n519_n5000#
+ a_n82_n5088# a_n225_n5000# a_363_n5000# a_408_5022# a_212_5022# a_n376_5022# a_n421_n5000#
+ a_n278_n5088# a_n127_n5000# a_265_n5000# a_n180_5022#
X0 a_n421_n5000# a_n474_n5088# a_n519_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X1 a_n225_n5000# a_n278_n5088# a_n323_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X2 a_69_n5000# a_16_5022# a_n29_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X3 a_167_n5000# a_114_n5088# a_69_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=0p ps=0u w=5e+07u l=200000u
X4 a_363_n5000# a_310_n5088# a_265_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X5 a_n29_n5000# a_n82_n5088# a_n127_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X6 a_n323_n5000# a_n376_5022# a_n421_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X7 a_n127_n5000# a_n180_5022# a_n225_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X8 a_265_n5000# a_212_5022# a_167_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X9 a_461_n5000# a_408_5022# a_363_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=0p ps=0u w=5e+07u l=200000u
.ends

.subckt diode_connected_nmos m1_60_4610# m1_120_80# VSUBS
Xsky130_fd_pr__nfet_01v8_UXPKRJ_0 VSUBS m1_120_80# m1_120_80# m1_120_80# m1_60_4610#
+ m1_60_4610# m1_120_80# m1_60_4610# m1_120_80# m1_120_80# m1_60_4610# m1_120_80#
+ m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_60_4610#
+ m1_60_4610# m1_120_80# sky130_fd_pr__nfet_01v8_UXPKRJ
.ends

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VPWR Y VNB VPB
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=2.05e+12p pd=1.41e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_BDZ9JN a_15_n500# a_n177_n500# a_n561_n500# a_879_n500#
+ a_111_n500# a_n129_n597# a_n513_n597# a_n609_531# a_63_n597# a_n273_n500# a_n801_531#
+ a_687_n500# a_n321_n597# a_159_531# a_639_n597# a_n941_n500# a_783_n500# a_399_n500#
+ a_n81_n500# a_n849_n500# a_351_531# a_n33_531# a_495_n500# a_n897_n597# a_831_n597#
+ a_447_n597# a_n225_531# a_591_n500# a_n657_n500# a_207_n500# a_543_531# a_n753_n500#
+ a_n369_n500# a_303_n500# a_255_n597# a_n705_n597# a_n417_531# w_n1079_n719# a_n465_n500#
+ a_735_531#
X0 a_15_n500# a_n33_531# a_n81_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X1 a_n369_n500# a_n417_531# a_n465_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X2 a_n657_n500# a_n705_n597# a_n753_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X3 a_879_n500# a_831_n597# a_783_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.55e+12p pd=1.062e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X4 a_303_n500# a_255_n597# a_207_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X5 a_n273_n500# a_n321_n597# a_n369_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X6 a_591_n500# a_543_531# a_495_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X7 a_n849_n500# a_n897_n597# a_n941_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.55e+12p ps=1.062e+07u w=5e+06u l=150000u
X8 a_207_n500# a_159_531# a_111_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X9 a_n177_n500# a_n225_531# a_n273_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X10 a_495_n500# a_447_n597# a_399_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X11 a_n561_n500# a_n609_531# a_n657_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X12 a_111_n500# a_63_n597# a_15_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X13 a_783_n500# a_735_531# a_687_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X14 a_399_n500# a_351_531# a_303_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X15 a_n465_n500# a_n513_n597# a_n561_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X16 a_687_n500# a_639_n597# a_591_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X17 a_n753_n500# a_n801_531# a_n849_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X18 a_n81_n500# a_n129_n597# a_n177_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_KBNS5F a_15_n500# a_n177_n500# a_111_n500# a_n273_n500#
+ a_159_n588# a_63_522# a_255_522# a_399_n500# a_n81_n500# a_351_n588# a_n417_n588#
+ a_n129_522# a_n225_n588# a_n321_522# a_n563_n674# a_207_n500# a_n461_n500# a_n369_n500#
+ a_303_n500# a_n33_n588#
X0 a_n81_n500# a_n129_522# a_n177_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X1 a_15_n500# a_n33_n588# a_n81_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X2 a_n369_n500# a_n417_n588# a_n461_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.55e+12p ps=1.062e+07u w=5e+06u l=150000u
X3 a_n273_n500# a_n321_522# a_n369_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X4 a_303_n500# a_255_522# a_207_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X5 a_n177_n500# a_n225_n588# a_n273_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6 a_207_n500# a_159_n588# a_111_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X7 a_111_n500# a_63_522# a_15_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8 a_399_n500# a_351_n588# a_303_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.55e+12p pd=1.062e+07u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sized_switch m1_970_n860# m1_1100_n50# m1_1190_n720# m1_3210_n860# w_2760_n990#
+ VSUBS
XXM1 m1_1100_n50# m1_1100_n50# m1_1100_n50# m1_1190_n720# m1_1190_n720# m1_970_n860#
+ m1_970_n860# m1_970_n860# m1_970_n860# m1_1190_n720# m1_970_n860# m1_1190_n720#
+ m1_970_n860# m1_970_n860# m1_970_n860# m1_1100_n50# m1_1100_n50# m1_1100_n50# m1_1190_n720#
+ m1_1190_n720# m1_970_n860# m1_970_n860# m1_1190_n720# m1_970_n860# m1_970_n860#
+ m1_970_n860# m1_970_n860# m1_1100_n50# m1_1190_n720# m1_1100_n50# m1_970_n860# m1_1100_n50#
+ m1_1100_n50# m1_1190_n720# m1_970_n860# m1_970_n860# m1_970_n860# w_2760_n990# m1_1190_n720#
+ m1_970_n860# sky130_fd_pr__pfet_01v8_BDZ9JN
Xsky130_fd_pr__nfet_01v8_KBNS5F_0 m1_1190_n720# m1_1190_n720# m1_1100_n50# m1_1100_n50#
+ m1_3210_n860# m1_3210_n860# m1_3210_n860# m1_1190_n720# m1_1100_n50# m1_3210_n860#
+ m1_3210_n860# m1_3210_n860# m1_3210_n860# m1_3210_n860# VSUBS m1_1190_n720# m1_1100_n50#
+ m1_1190_n720# m1_1100_n50# m1_3210_n860# sky130_fd_pr__nfet_01v8_KBNS5F
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt analog_mux OUT VDD SIG0 SIG1 SIG2 SIG3 SIG4 SIG5 SIG6 SIG7 SIG8 SIG9 SIG10
+ SIG11 SIG12 SIG13 SIG14 SIG15 SEL0 SEL1 SEL2 SEL3 GND
Xx1 x8/A x9/B x9/C x9/D GND VDD x1/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx2 x8/A x9/B x9/C SEL0 GND VDD x2/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx3 x8/A x9/B SEL1 x9/D GND VDD x3/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx4 x8/A x9/B SEL1 SEL0 GND VDD x4/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx5 x8/A SEL2 x9/C x9/D GND VDD x5/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx6 x8/A SEL2 x9/C SEL0 GND VDD x6/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_0 x7/Y OUT SIG6 sky130_fd_sc_hd__inv_2_15/Y VDD GND sized_switch
Xsized_switch_1 x2/Y OUT SIG1 sky130_fd_sc_hd__inv_2_2/Y VDD GND sized_switch
Xx7 x8/A SEL2 SEL1 x9/D GND VDD x7/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_2 x3/Y OUT SIG2 sky130_fd_sc_hd__inv_2_3/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_10 x12/Y GND VDD sky130_fd_sc_hd__inv_2_10/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_11 x13/Y GND VDD sky130_fd_sc_hd__inv_2_11/Y GND VDD sky130_fd_sc_hd__inv_2
Xx8 x8/A SEL2 SEL1 SEL0 GND VDD x8/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_3 x4/Y OUT SIG3 sky130_fd_sc_hd__inv_2_0/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_12 x14/Y GND VDD sky130_fd_sc_hd__inv_2_12/Y GND VDD sky130_fd_sc_hd__inv_2
Xx9 SEL3 x9/B x9/C x9/D GND VDD x9/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_4 x5/Y OUT SIG4 sky130_fd_sc_hd__inv_2_5/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_13 x15/Y GND VDD sky130_fd_sc_hd__inv_2_13/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_5 x6/Y OUT SIG5 sky130_fd_sc_hd__inv_2_6/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_14 x16/Y GND VDD sky130_fd_sc_hd__inv_2_14/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_6 x11/Y OUT SIG10 sky130_fd_sc_hd__inv_2_9/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_0 x4/Y GND VDD sky130_fd_sc_hd__inv_2_0/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_15 x7/Y GND VDD sky130_fd_sc_hd__inv_2_15/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_7 x10/Y OUT SIG9 sky130_fd_sc_hd__inv_2_8/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_1 x8/Y GND VDD sky130_fd_sc_hd__inv_2_1/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_8 x12/Y OUT SIG11 sky130_fd_sc_hd__inv_2_10/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_2 x2/Y GND VDD sky130_fd_sc_hd__inv_2_2/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_9 x13/Y OUT SIG12 sky130_fd_sc_hd__inv_2_11/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_3 x3/Y GND VDD sky130_fd_sc_hd__inv_2_3/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_4 x1/Y GND VDD sky130_fd_sc_hd__inv_2_4/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_5 x5/Y GND VDD sky130_fd_sc_hd__inv_2_5/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_6 x6/Y GND VDD sky130_fd_sc_hd__inv_2_6/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_7 x9/Y GND VDD sky130_fd_sc_hd__inv_2_7/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_8 x10/Y GND VDD sky130_fd_sc_hd__inv_2_8/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_9 x11/Y GND VDD sky130_fd_sc_hd__inv_2_9/Y GND VDD sky130_fd_sc_hd__inv_2
Xx20 SEL0 GND VDD x9/D GND VDD sky130_fd_sc_hd__inv_8
Xx10 SEL3 x9/B x9/C SEL0 GND VDD x10/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_10 x14/Y OUT SIG13 sky130_fd_sc_hd__inv_2_12/Y VDD GND sized_switch
Xx11 SEL3 x9/B SEL1 x9/D GND VDD x11/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_11 x15/Y OUT SIG14 sky130_fd_sc_hd__inv_2_13/Y VDD GND sized_switch
Xx12 SEL3 x9/B SEL1 SEL0 GND VDD x12/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_12 x8/Y OUT SIG7 sky130_fd_sc_hd__inv_2_1/Y VDD GND sized_switch
Xx13 SEL3 SEL2 x9/C x9/D GND VDD x13/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_13 x9/Y OUT SIG8 sky130_fd_sc_hd__inv_2_7/Y VDD GND sized_switch
Xx14 SEL3 SEL2 x9/C SEL0 GND VDD x14/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx15 SEL3 SEL2 SEL1 x9/D GND VDD x15/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_14 x1/Y OUT SIG0 sky130_fd_sc_hd__inv_2_4/Y VDD GND sized_switch
Xx16 SEL3 SEL2 SEL1 SEL0 GND VDD x16/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_15 x16/Y OUT SIG15 sky130_fd_sc_hd__inv_2_14/Y VDD GND sized_switch
Xx17 SEL3 GND VDD x8/A GND VDD sky130_fd_sc_hd__inv_8
Xx18 SEL2 GND VDD x9/B GND VDD sky130_fd_sc_hd__inv_8
Xx19 SEL1 GND VDD x9/C GND VDD sky130_fd_sc_hd__inv_8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_95KK7Z c1_n1650_n1600# m3_n1750_n1700#
X0 c1_n1650_n1600# m3_n1750_n1700# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_49C6SK a_n50_n596# a_524_n500# a_n682_n596# a_1214_n596#
+ a_n1472_n596# a_1156_n500# a_740_n596# a_682_n500# a_50_n500# a_1372_n596# a_n840_n596#
+ a_n1630_n596# a_1314_n500# a_840_n500# a_n108_n500# a_1530_n596# a_1472_n500# a_n266_n500#
+ a_n898_n500# a_n1056_n500# a_1630_n500# a_n1688_n500# a_108_n596# a_n424_n500# a_n208_n596#
+ a_n1214_n500# w_n1826_n718# a_n582_n500# a_266_n596# a_208_n500# a_n1372_n500# a_898_n596#
+ a_n366_n596# a_424_n596# a_n998_n596# a_n1156_n596# a_n740_n500# a_366_n500# a_n1530_n500#
+ a_1056_n596# a_n524_n596# a_998_n500# a_582_n596# a_n1314_n596#
X0 a_524_n500# a_424_n596# a_366_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_1630_n500# a_1530_n596# a_1472_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_n1056_n500# a_n1156_n596# a_n1214_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_1156_n500# a_1056_n596# a_998_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_n108_n500# a_n208_n596# a_n266_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_208_n500# a_108_n596# a_50_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1214_n500# a_n1314_n596# a_n1372_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1314_n500# a_1214_n596# a_1156_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X8 a_n740_n500# a_n840_n596# a_n898_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_n582_n500# a_n682_n596# a_n740_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X10 a_682_n500# a_582_n596# a_524_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n266_n500# a_n366_n596# a_n424_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_840_n500# a_740_n596# a_682_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n1530_n500# a_n1630_n596# a_n1688_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_366_n500# a_266_n596# a_208_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_n1372_n500# a_n1472_n596# a_n1530_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_1472_n500# a_1372_n596# a_1314_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_n898_n500# a_n998_n596# a_n1056_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_50_n500# a_n50_n596# a_n108_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_n424_n500# a_n524_n596# a_n582_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 a_998_n500# a_898_n596# a_840_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_JT3SH9 a_n1318_n500# a_1060_n588# a_n286_n500# a_n1060_n500#
+ a_n1518_n588# a_n486_n588# a_744_n500# a_n1260_n588# a_544_n588# a_1776_n500# a_1576_n588#
+ a_228_n500# a_n1576_n500# a_n544_n500# a_28_n588# a_n1776_n588# a_n744_n588# a_1002_n500#
+ a_802_n588# a_n1936_n674# a_486_n500# a_n28_n500# a_n228_n588# a_n1834_n500# a_286_n588#
+ a_n1002_n588# a_1518_n500# a_n802_n500# a_1260_n500# a_1318_n588#
X0 a_n1318_n500# a_n1518_n588# a_n1576_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_n544_n500# a_n744_n588# a_n802_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_n1060_n500# a_n1260_n588# a_n1318_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X3 a_n286_n500# a_n486_n588# a_n544_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X4 a_n802_n500# a_n1002_n588# a_n1060_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 a_n1576_n500# a_n1776_n588# a_n1834_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X6 a_1518_n500# a_1318_n588# a_1260_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X7 a_1002_n500# a_802_n588# a_744_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X8 a_486_n500# a_286_n588# a_228_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X9 a_744_n500# a_544_n588# a_486_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X10 a_1776_n500# a_1576_n588# a_1518_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X11 a_1260_n500# a_1060_n588# a_1002_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 a_228_n500# a_28_n588# a_n28_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.4e+12p ps=1.056e+07u w=5e+06u l=1e+06u
X13 a_n28_n500# a_n228_n588# a_n286_n500# a_n1936_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_F7BMVG a_n573_n1432# a_n703_n1562# a_n573_1000#
X0 a_n573_n1432# a_n573_1000# a_n703_n1562# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_JEXVB9 a_1261_n500# a_1319_n588# a_n1319_n500# a_1061_n588#
+ a_n287_n500# a_n1061_n500# a_n1519_n588# a_n487_n588# a_745_n500# a_n1261_n588#
+ a_545_n588# a_n1679_n674# a_229_n500# a_n1577_n500# a_n545_n500# a_29_n588# a_1003_n500#
+ a_n745_n588# a_803_n588# a_n29_n500# a_487_n500# a_n229_n588# a_n1003_n588# a_287_n588#
+ a_1519_n500# a_n803_n500#
X0 a_1519_n500# a_1319_n588# a_1261_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_n1061_n500# a_n1261_n588# a_n1319_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_1003_n500# a_803_n588# a_745_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_487_n500# a_287_n588# a_229_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_745_n500# a_545_n588# a_487_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 a_1261_n500# a_1061_n588# a_1003_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 a_n29_n500# a_n229_n588# a_n287_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X7 a_229_n500# a_29_n588# a_n29_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 a_n1319_n500# a_n1519_n588# a_n1577_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X9 a_n545_n500# a_n745_n588# a_n803_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X10 a_n803_n500# a_n1003_n588# a_n1061_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X11 a_n287_n500# a_n487_n588# a_n545_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_EJ3ASN a_524_n500# a_108_n588# a_50_n500# a_n208_n588#
+ a_266_n588# a_n366_n588# a_n108_n500# a_424_n588# a_n524_n588# a_n266_n500# a_n50_n588#
+ a_n424_n500# a_n684_n674# a_n582_n500# a_208_n500# a_366_n500#
X0 a_366_n500# a_266_n588# a_208_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n500# a_n50_n588# a_n108_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_n424_n500# a_n524_n588# a_n582_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_524_n500# a_424_n588# a_366_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X4 a_n108_n500# a_n208_n588# a_n266_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_208_n500# a_108_n588# a_50_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X6 a_n266_n500# a_n366_n588# a_n424_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_9F67JW a_n1608_n500# a_28_n596# a_n976_n500# a_n1134_n500#
+ a_n128_n596# a_n2556_n500# a_186_n596# a_n1766_n500# a_n2082_n500# a_128_n500# a_n502_n500#
+ a_n1292_n500# a_818_n596# a_n286_n596# a_n1076_n596# a_n2714_n500# a_n3030_n500#
+ a_344_n596# a_n2498_n596# a_286_n500# a_n660_n500# a_n1924_n500# a_n2240_n500# a_n918_n596#
+ a_976_n596# a_n444_n596# a_n1450_n500# a_n1708_n596# a_n2024_n596# a_n2872_n500#
+ a_2398_n596# a_n1234_n596# a_918_n500# a_502_n596# a_n2656_n596# a_444_n500# a_1608_n596#
+ a_n1866_n596# a_n602_n596# a_n2182_n596# a_1134_n596# a_660_n596# a_n1392_n596#
+ a_1076_n500# a_2556_n596# a_2498_n500# a_2082_n596# a_1766_n596# a_n2814_n596# a_602_n500#
+ a_1292_n596# a_n760_n596# a_n3130_n596# a_1708_n500# a_n2340_n596# a_2024_n500#
+ a_n1550_n596# a_1234_n500# a_3030_n596# a_2714_n596# a_n2972_n596# a_2656_n500#
+ a_760_n500# a_2240_n596# a_1924_n596# a_2182_n500# a_1866_n500# a_1450_n596# a_1392_n500#
+ a_n28_n500# a_2872_n596# a_n186_n500# a_3130_n500# a_2814_n500# a_2340_n500# a_n3188_n500#
+ a_1550_n500# a_n2398_n500# a_2972_n500# a_n818_n500# a_n344_n500# w_n3326_n718#
X0 a_n1134_n500# a_n1234_n596# a_n1292_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n660_n500# a_n760_n596# a_n818_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_1234_n500# a_1134_n596# a_1076_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n2714_n500# a_n2814_n596# a_n2872_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_2814_n500# a_2714_n596# a_2656_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_3130_n500# a_3030_n596# a_2972_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n2240_n500# a_n2340_n596# a_n2398_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_n1766_n500# a_n1866_n596# a_n1924_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_1866_n500# a_1766_n596# a_1708_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_n2082_n500# a_n2182_n596# a_n2240_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X10 a_2182_n500# a_2082_n596# a_2024_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X11 a_n818_n500# a_n918_n596# a_n976_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_918_n500# a_818_n596# a_760_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X13 a_n186_n500# a_n286_n596# a_n344_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_760_n500# a_660_n596# a_602_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X15 a_2024_n500# a_1924_n596# a_1866_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_2340_n500# a_2240_n596# a_2182_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X17 a_n1450_n500# a_n1550_n596# a_n1608_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X18 a_286_n500# a_186_n596# a_128_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X19 a_n1292_n500# a_n1392_n596# a_n1450_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 a_1392_n500# a_1292_n596# a_1234_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X21 a_n2872_n500# a_n2972_n596# a_n3030_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X22 a_2972_n500# a_2872_n596# a_2814_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X23 a_n344_n500# a_n444_n596# a_n502_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X24 a_n2398_n500# a_n2498_n596# a_n2556_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X25 a_2498_n500# a_2398_n596# a_2340_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X26 a_128_n500# a_28_n596# a_n28_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.4e+12p ps=1.056e+07u w=5e+06u l=500000u
X27 a_n1608_n500# a_n1708_n596# a_n1766_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X28 a_444_n500# a_344_n596# a_286_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X29 a_1708_n500# a_1608_n596# a_1550_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X30 a_n1924_n500# a_n2024_n596# a_n2082_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X31 a_1550_n500# a_1450_n596# a_1392_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X32 a_n976_n500# a_n1076_n596# a_n1134_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X33 a_1076_n500# a_976_n596# a_918_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X34 a_n3030_n500# a_n3130_n596# a_n3188_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X35 a_n2556_n500# a_n2656_n596# a_n2714_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X36 a_n502_n500# a_n602_n596# a_n660_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X37 a_2656_n500# a_2556_n596# a_2498_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X38 a_n28_n500# a_n128_n596# a_n186_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X39 a_602_n500# a_502_n596# a_444_n500# w_n3326_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_GNAJ57 a_n50_n596# a_524_n500# a_n682_n596# a_1214_n596#
+ a_n1472_n596# a_1156_n500# a_740_n596# a_682_n500# a_50_n500# a_1372_n596# a_n840_n596#
+ a_n1630_n596# a_1314_n500# a_840_n500# a_n108_n500# a_1530_n596# a_1472_n500# a_n266_n500#
+ a_n898_n500# a_n1056_n500# a_1630_n500# a_n1688_n500# a_108_n596# a_n424_n500# a_n208_n596#
+ a_n1214_n500# w_n1826_n718# a_n582_n500# a_266_n596# a_208_n500# a_n1372_n500# a_898_n596#
+ a_n366_n596# a_424_n596# a_n998_n596# a_n1156_n596# a_n740_n500# a_366_n500# a_n1530_n500#
+ a_1056_n596# a_n524_n596# a_998_n500# a_582_n596# a_n1314_n596#
X0 a_524_n500# a_424_n596# a_366_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_1630_n500# a_1530_n596# a_1472_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_n1056_n500# a_n1156_n596# a_n1214_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_1156_n500# a_1056_n596# a_998_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_n108_n500# a_n208_n596# a_n266_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_208_n500# a_108_n596# a_50_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1214_n500# a_n1314_n596# a_n1372_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1314_n500# a_1214_n596# a_1156_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X8 a_n740_n500# a_n840_n596# a_n898_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_n582_n500# a_n682_n596# a_n740_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X10 a_682_n500# a_582_n596# a_524_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n266_n500# a_n366_n596# a_n424_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_840_n500# a_740_n596# a_682_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n1530_n500# a_n1630_n596# a_n1688_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_366_n500# a_266_n596# a_208_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_n1372_n500# a_n1472_n596# a_n1530_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_1472_n500# a_1372_n596# a_1314_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_n898_n500# a_n998_n596# a_n1056_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_50_n500# a_n50_n596# a_n108_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_n424_n500# a_n524_n596# a_n582_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 a_998_n500# a_898_n596# a_840_n500# w_n1826_n718# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt OTA_fingers_031123_NON_FLAT m1_n1130_9530# m1_1130_3110# li_900_7430# m1_n500_70#
+ m1_1130_4630# VSUBS
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_2 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_3 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__pfet_01v8_49C6SK_0 m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730#
+ m1_90_7730# li_900_7430# m1_90_7730# m1_n2620_8810# m1_n2620_8810# m1_90_7730# m1_90_7730#
+ m1_90_7730# m1_n2620_8810# li_900_7430# li_900_7430# m1_90_7730# li_900_7430# m1_n2620_8810#
+ m1_n2620_8810# li_900_7430# m1_n2620_8810# li_900_7430# m1_90_7730# li_900_7430#
+ m1_90_7730# m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_90_7730# li_900_7430#
+ li_900_7430# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# li_900_7430#
+ m1_n2620_8810# m1_n2620_8810# m1_90_7730# m1_90_7730# m1_n2620_8810# m1_90_7730#
+ m1_90_7730# sky130_fd_pr__pfet_01v8_49C6SK
Xsky130_fd_pr__nfet_01v8_JT3SH9_0 m1_60_860# m1_n500_70# m1_60_860# VSUBS m1_n500_70#
+ m1_n500_70# m1_60_860# m1_n500_70# m1_n500_70# m1_60_860# m1_n500_70# m1_60_860#
+ VSUBS VSUBS m1_n500_70# m1_n500_70# m1_n500_70# VSUBS m1_n500_70# VSUBS VSUBS VSUBS
+ m1_n500_70# m1_60_860# m1_n500_70# m1_n500_70# VSUBS m1_60_860# m1_60_860# m1_n500_70#
+ sky130_fd_pr__nfet_01v8_JT3SH9
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0 m1_n5940_10010# VSUBS m1_n2620_8810# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1 m1_n5940_10010# VSUBS m1_n2620_8810# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2 m1_n2620_8810# VSUBS m1_n5940_10010# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__nfet_01v8_JEXVB9_0 VSUBS m1_n500_70# VSUBS m1_n500_70# VSUBS m1_n1130_9530#
+ m1_n500_70# m1_n500_70# VSUBS m1_n500_70# m1_n500_70# VSUBS VSUBS m1_n1130_9530#
+ m1_n1130_9530# m1_n500_70# m1_n1130_9530# m1_n500_70# m1_n500_70# m1_n1130_9530#
+ m1_n1130_9530# m1_n500_70# m1_n500_70# m1_n500_70# m1_n1130_9530# VSUBS sky130_fd_pr__nfet_01v8_JEXVB9
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3 m1_n2620_8810# VSUBS m1_n5940_10010# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__nfet_01v8_EJ3ASN_0 m1_60_860# m1_1130_4630# m1_n2620_8810# m1_1130_4630#
+ m1_1130_4630# m1_1130_4630# m1_60_860# m1_1130_4630# m1_1130_4630# m1_n2620_8810#
+ m1_1130_4630# m1_60_860# VSUBS m1_n2620_8810# m1_60_860# m1_n2620_8810# sky130_fd_pr__nfet_01v8_EJ3ASN
Xsky130_fd_pr__pfet_01v8_9F67JW_0 li_900_7430# m1_n2620_8810# li_900_7430# m1_n1130_9530#
+ m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_n1130_9530# m1_n1130_9530# m1_n1130_9530#
+ m1_n1130_9530# li_900_7430# m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_n1130_9530#
+ m1_n1130_9530# m1_n2620_8810# m1_n2620_8810# li_900_7430# li_900_7430# li_900_7430#
+ li_900_7430# m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_n1130_9530# m1_n2620_8810#
+ m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_n2620_8810# li_900_7430# m1_n2620_8810#
+ m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_n2620_8810#
+ m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# li_900_7430#
+ m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_n2620_8810#
+ m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# li_900_7430#
+ m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_n1130_9530# m1_n1130_9530# m1_n2620_8810#
+ m1_n2620_8810# li_900_7430# li_900_7430# m1_n2620_8810# m1_n1130_9530# li_900_7430#
+ m1_n2620_8810# m1_n1130_9530# li_900_7430# li_900_7430# m1_n1130_9530# li_900_7430#
+ li_900_7430# m1_n1130_9530# m1_n1130_9530# m1_n1130_9530# li_900_7430# li_900_7430#
+ sky130_fd_pr__pfet_01v8_9F67JW
Xsky130_fd_pr__nfet_01v8_EJ3ASN_1 m1_90_7730# m1_1130_3110# m1_60_860# m1_1130_3110#
+ m1_1130_3110# m1_1130_3110# m1_90_7730# m1_1130_3110# m1_1130_3110# m1_60_860# m1_1130_3110#
+ m1_90_7730# VSUBS m1_60_860# m1_90_7730# m1_60_860# sky130_fd_pr__nfet_01v8_EJ3ASN
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_0 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__pfet_01v8_GNAJ57_0 m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730#
+ m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730#
+ m1_90_7730# m1_90_7730# li_900_7430# li_900_7430# m1_90_7730# li_900_7430# m1_90_7730#
+ m1_90_7730# li_900_7430# m1_90_7730# li_900_7430# m1_90_7730# li_900_7430# m1_90_7730#
+ m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730# li_900_7430# li_900_7430# m1_90_7730#
+ m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730#
+ m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# sky130_fd_pr__pfet_01v8_GNAJ57
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_1 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
.ends

.subckt constant_gm_local_030423 a_n3719_36# w_n4170_1941# a_n3633_196#
X0 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X1 a_n3688_2136# a_n3688_2136# a_n3633_196# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.348e+07u w=2.5e+06u l=500000u
X2 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=1.74e+13p pd=1.2696e+08u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X3 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X5 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.232e+07u w=1.25e+06u l=1e+06u
X6 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X7 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X9 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X10 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X11 a_n3688_2136# a_n3688_2136# a_n3633_196# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X12 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X14 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X17 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X20 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X21 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X22 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X23 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X24 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X25 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X26 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X27 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_SDAUVS a_n50_n2451# a_n108_n2354# a_n108_118# a_n108_1354#
+ a_n50_1257# a_n50_21# a_n50_4965# a_50_3826# a_50_118# a_50_n3590# a_n50_n1215#
+ a_50_n6062# a_n50_n4923# a_n108_n1118# a_n108_3826# w_n246_n6281# a_n108_n4826#
+ a_n50_n3687# a_n50_3729# a_n50_n6159# a_50_2590# a_50_n2354# a_50_5062# a_n108_2590#
+ a_n108_n3590# a_n50_2493# a_n108_5062# a_n108_n6062# a_50_1354# a_50_n1118# a_50_n4826#
X0 a_50_n6062# a_n50_n6159# a_n108_n6062# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_2590# a_n50_2493# a_n108_2590# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_118# a_n50_21# a_n108_118# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_5062# a_n50_4965# a_n108_5062# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_n4826# a_n50_n4923# a_n108_n4826# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_n2354# a_n50_n2451# a_n108_n2354# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_3826# a_n50_3729# a_n108_3826# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_50_1354# a_n50_1257# a_n108_1354# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_50_n1118# a_n50_n1215# a_n108_n1118# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_50_n3590# a_n50_n3687# a_n108_n3590# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_K6FQWW a_n108_1936# a_n108_n2936# a_n108_718# a_50_n500#
+ a_n50_n3024# a_50_3154# a_n210_n4328# a_50_718# a_n108_n500# a_n50_630# a_n108_n1718#
+ a_n108_3154# a_n108_n4154# a_n50_n588# a_50_n2936# a_n50_1848# a_n50_n1806# a_n50_n4242#
+ a_50_1936# a_50_n1718# a_50_n4154# a_n50_3066#
X0 a_50_n2936# a_n50_n3024# a_n108_n2936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n500# a_n50_n588# a_n108_n500# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_n4154# a_n50_n4242# a_n108_n4154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_1936# a_n50_1848# a_n108_1936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_3154# a_n50_3066# a_n108_3154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_718# a_n50_630# a_n108_718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_n1718# a_n50_n1806# a_n108_n1718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_KG6QWW a_n100_3066# a_n158_1936# a_100_n1718# a_100_n4154#
+ a_100_n500# a_n100_n3024# a_n158_718# a_100_3154# a_n158_n2936# a_n158_n500# a_n158_3154#
+ a_n260_n4328# a_n100_n588# a_n158_n1718# a_n100_1848# a_n158_n4154# a_100_718# a_n100_630#
+ a_100_n2936# a_n100_n4242# a_n100_n1806# a_100_1936#
X0 a_100_718# a_n100_630# a_n158_718# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_100_1936# a_n100_1848# a_n158_1936# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_100_n1718# a_n100_n1806# a_n158_n1718# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_100_3154# a_n100_3066# a_n158_3154# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_100_n2936# a_n100_n3024# a_n158_n2936# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X6 a_100_n4154# a_n100_n4242# a_n158_n4154# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_T9YF2H a_n50_n597# w_n246_n4427# a_n108_n2972# a_50_n500#
+ a_n108_736# a_n108_1972# a_n50_1875# a_50_3208# a_n108_n500# a_50_736# a_n50_n1833#
+ a_n50_n4305# a_n108_n1736# a_n108_n4208# a_n50_n3069# a_n108_3208# a_n50_639# a_50_n2972#
+ a_n50_3111# a_50_1972# a_50_n1736# a_50_n4208#
X0 a_50_736# a_n50_639# a_n108_736# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n2972# a_n50_n3069# a_n108_n2972# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_1972# a_n50_1875# a_n108_1972# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_n1736# a_n50_n1833# a_n108_n1736# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_n4208# a_n50_n4305# a_n108_n4208# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_3208# a_n50_3111# a_n108_3208# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_n500# a_n50_n597# a_n108_n500# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_GG6QWW a_100_n3545# a_n100_n2415# a_100_2545# a_n100_n1197#
+ a_n158_n1109# a_n100_1239# a_n100_21# a_n260_n3719# a_100_109# a_n158_2545# a_100_n2327#
+ a_100_1327# a_n158_n3545# a_n158_1327# a_100_n1109# a_n100_n3633# a_n158_109# a_n158_n2327#
+ a_n100_2457#
X0 a_100_1327# a_n100_1239# a_n158_1327# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_100_2545# a_n100_2457# a_n158_2545# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_100_n1109# a_n100_n1197# a_n158_n1109# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_100_n2327# a_n100_n2415# a_n158_n2327# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_100_n3545# a_n100_n3633# a_n158_n3545# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_100_109# a_n100_21# a_n158_109# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_R8BLL7 a_n108_1936# a_n108_n2936# a_n108_718# a_50_n500#
+ a_n50_n3024# a_50_3154# a_n210_n4328# a_50_718# a_n108_n500# a_n50_630# a_n108_n1718#
+ a_n108_3154# a_n108_n4154# a_n50_n588# a_50_n2936# a_n50_1848# a_n50_n1806# a_n50_n4242#
+ a_50_1936# a_50_n1718# a_50_n4154# a_n50_3066#
X0 a_50_n2936# a_n50_n3024# a_n108_n2936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n500# a_n50_n588# a_n108_n500# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_n4154# a_n50_n4242# a_n108_n4154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_1936# a_n50_1848# a_n108_1936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_3154# a_n50_3066# a_n108_3154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_718# a_n50_630# a_n108_718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_n1718# a_n50_n1806# a_n108_n1718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt ota_3_11_23_nonflat m1_n6050_3760# m1_n4180_2590# m1_n4190_3090# m1_n4200_780#
+ w_n6280_3640# VSUBS
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_3 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_2 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__pfet_01v8_SDAUVS_0 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__pfet_01v8_SDAUVS_1 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__pfet_01v8_SDAUVS_2 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__pfet_01v8_SDAUVS_3 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__nfet_01v8_K6FQWW_0 m1_n4120_60# m1_n4120_60# m1_n4120_60# m1_n4300_8710#
+ m1_n4180_2590# m1_n4300_8710# VSUBS m1_n4300_8710# m1_n4120_60# m1_n4180_2590# m1_n4120_60#
+ m1_n4120_60# m1_n4120_60# m1_n4180_2590# m1_n4300_8710# m1_n4180_2590# m1_n4180_2590#
+ m1_n4180_2590# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4180_2590# sky130_fd_pr__nfet_01v8_K6FQWW
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0 m1_n7530_3520# VSUBS m1_n9960_3530# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1 m1_n7530_3520# VSUBS m1_n9960_3530# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__nfet_01v8_KG6QWW_0 m1_n4200_780# VSUBS m1_n4120_60# m1_n4120_60# m1_n4120_60#
+ m1_n4200_780# VSUBS m1_n4120_60# VSUBS VSUBS VSUBS VSUBS m1_n4200_780# VSUBS m1_n4200_780#
+ VSUBS m1_n4120_60# m1_n4200_780# m1_n4120_60# m1_n4200_780# m1_n4200_780# m1_n4120_60#
+ sky130_fd_pr__nfet_01v8_KG6QWW
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2 m1_n9960_3530# VSUBS m1_n7530_3520# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__nfet_01v8_KG6QWW_1 m1_n4200_780# VSUBS m1_n4120_60# m1_n4120_60# m1_n4120_60#
+ m1_n4200_780# VSUBS m1_n4120_60# VSUBS VSUBS VSUBS VSUBS m1_n4200_780# VSUBS m1_n4200_780#
+ VSUBS m1_n4120_60# m1_n4200_780# m1_n4120_60# m1_n4200_780# m1_n4200_780# m1_n4120_60#
+ sky130_fd_pr__nfet_01v8_KG6QWW
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3 m1_n9960_3530# VSUBS m1_n7530_3520# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__pfet_01v8_T9YF2H_0 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n7530_3520#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n7530_3520# w_n6280_3640# m1_n7530_3520#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n7530_3520# m1_n4300_8710# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_1 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n4300_8710# w_n6280_3640# m1_n4300_8710#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_2 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n7530_3520#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n7530_3520# w_n6280_3640# m1_n7530_3520#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n7530_3520# m1_n4300_8710# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_3 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n4300_8710# w_n6280_3640# m1_n4300_8710#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_5 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n7530_3520#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n7530_3520# w_n6280_3640# m1_n7530_3520#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n7530_3520# m1_n4300_8710# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_4 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n4300_8710# w_n6280_3640# m1_n4300_8710#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__nfet_01v8_GG6QWW_0 VSUBS m1_n4200_780# VSUBS m1_n4200_780# m1_n6050_3760#
+ m1_n4200_780# m1_n4200_780# VSUBS VSUBS m1_n6050_3760# VSUBS VSUBS m1_n6050_3760#
+ m1_n6050_3760# VSUBS m1_n4200_780# m1_n6050_3760# m1_n6050_3760# m1_n4200_780# sky130_fd_pr__nfet_01v8_GG6QWW
Xsky130_fd_pr__nfet_01v8_R8BLL7_0 m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n4120_60#
+ m1_n4190_3090# m1_n4120_60# VSUBS m1_n4120_60# m1_n7530_3520# m1_n4190_3090# m1_n7530_3520#
+ m1_n7530_3520# m1_n7530_3520# m1_n4190_3090# m1_n4120_60# m1_n4190_3090# m1_n4190_3090#
+ m1_n4190_3090# m1_n4120_60# m1_n4120_60# m1_n4120_60# m1_n4190_3090# sky130_fd_pr__nfet_01v8_R8BLL7
Xsky130_fd_pr__nfet_01v8_GG6QWW_1 VSUBS m1_n4200_780# VSUBS m1_n4200_780# m1_n6050_3760#
+ m1_n4200_780# m1_n4200_780# VSUBS VSUBS m1_n6050_3760# VSUBS VSUBS m1_n6050_3760#
+ m1_n6050_3760# VSUBS m1_n4200_780# m1_n6050_3760# m1_n6050_3760# m1_n4200_780# sky130_fd_pr__nfet_01v8_GG6QWW
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_0 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_1 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
.ends

.subckt OTA_MULT_GM ota_3_11_23_nonflat_0/w_n6280_3640# ota_3_11_23_nonflat_0/m1_n4180_2590#
+ ota_3_11_23_nonflat_0/m1_n4190_3090# constant_gm_local_030423_0/w_n4170_1941# ota_3_11_23_nonflat_0/m1_n6050_3760#
+ VSUBS
Xconstant_gm_local_030423_0 VSUBS constant_gm_local_030423_0/w_n4170_1941# m1_n200_1910#
+ constant_gm_local_030423
Xota_3_11_23_nonflat_0 ota_3_11_23_nonflat_0/m1_n6050_3760# ota_3_11_23_nonflat_0/m1_n4180_2590#
+ ota_3_11_23_nonflat_0/m1_n4190_3090# m1_n200_1910# ota_3_11_23_nonflat_0/w_n6280_3640#
+ VSUBS ota_3_11_23_nonflat
.ends

.subckt sky130_fd_pr__nfet_01v8_A5635U a_n544_n124# a_n486_n212# a_486_n124# a_n28_n124#
+ a_28_n212# a_n286_n124# a_n228_n212# a_286_n212# a_228_n124# a_n646_n298#
X0 a_n286_n124# a_n486_n212# a_n544_n124# a_n646_n298# sky130_fd_pr__nfet_01v8 ad=3.596e+11p pd=3.06e+06u as=3.596e+11p ps=3.06e+06u w=1.24e+06u l=1e+06u
X1 a_486_n124# a_286_n212# a_228_n124# a_n646_n298# sky130_fd_pr__nfet_01v8 ad=3.596e+11p pd=3.06e+06u as=3.596e+11p ps=3.06e+06u w=1.24e+06u l=1e+06u
X2 a_228_n124# a_28_n212# a_n28_n124# a_n646_n298# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.472e+11p ps=3.04e+06u w=1.24e+06u l=1e+06u
X3 a_n28_n124# a_n228_n212# a_n286_n124# a_n646_n298# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_H7FLKU a_n28_n250# a_28_n338# a_n128_n338# a_n186_n250#
+ a_n288_n424# a_128_n250#
X0 a_n28_n250# a_n128_n338# a_n186_n250# a_n288_n424# sky130_fd_pr__nfet_01v8 ad=7e+11p pd=5.56e+06u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=500000u
X1 a_128_n250# a_28_n338# a_n28_n250# a_n288_n424# sky130_fd_pr__nfet_01v8 ad=7.25e+11p pd=5.58e+06u as=0p ps=0u w=2.5e+06u l=500000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_B5N4SD a_n572_6900# a_n572_n7332# VSUBS
X0 a_n572_n7332# a_n572_6900# VSUBS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_LK874N a_29_n597# a_n287_n500# a_n745_n597# a_745_n500#
+ a_n229_n597# a_287_n597# a_229_n500# a_n545_n500# w_n941_n719# a_n487_n597# a_n29_n500#
+ a_545_n597# a_487_n500# a_n803_n500#
X0 a_n29_n500# a_n229_n597# a_n287_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_229_n500# a_29_n597# a_n29_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X2 a_n545_n500# a_n745_n597# a_n803_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_n287_n500# a_n487_n597# a_n545_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 a_745_n500# a_545_n597# a_487_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_487_n500# a_287_n597# a_229_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_GLZPWL a_n286_n500# a_n486_n588# a_744_n500# a_544_n588#
+ a_228_n500# a_n544_n500# a_28_n588# a_n744_n588# a_486_n500# a_n28_n500# a_n228_n588#
+ a_286_n588# a_n904_n674# a_n802_n500#
X0 a_n544_n500# a_n744_n588# a_n802_n500# a_n904_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_n286_n500# a_n486_n588# a_n544_n500# a_n904_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X2 a_486_n500# a_286_n588# a_228_n500# a_n904_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_744_n500# a_544_n588# a_486_n500# a_n904_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X4 a_228_n500# a_28_n588# a_n28_n500# a_n904_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.4e+12p ps=1.056e+07u w=5e+06u l=1e+06u
X5 a_n28_n500# a_n228_n588# a_n286_n500# a_n904_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt constant_gm_fingers Vout VDD VSS
Xsky130_fd_pr__nfet_01v8_A5635U_0 VSS Vout VSS VSS Vout Vout Vout Vout Vout VSS sky130_fd_pr__nfet_01v8_A5635U
Xsky130_fd_pr__nfet_01v8_H7FLKU_0 Vout m1_n210_n170# m1_n210_n170# m1_n210_n170# VSS
+ m1_n210_n170# sky130_fd_pr__nfet_01v8_H7FLKU
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_0 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_1 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_2 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_3 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__pfet_01v8_LK874N_0 m1_n210_n170# VDD m1_n210_n170# VDD m1_n210_n170#
+ m1_n210_n170# VDD Vout VDD m1_n210_n170# Vout m1_n210_n170# Vout VDD sky130_fd_pr__pfet_01v8_LK874N
Xsky130_fd_pr__pfet_01v8_LK874N_1 m1_n210_n170# VDD m1_n210_n170# VDD m1_n210_n170#
+ m1_n210_n170# VDD m1_n210_n170# VDD m1_n210_n170# m1_n210_n170# m1_n210_n170# m1_n210_n170#
+ VDD sky130_fd_pr__pfet_01v8_LK874N
Xsky130_fd_pr__nfet_01v8_GLZPWL_0 m1_n210_n170# Vout m1_n210_n170# Vout m1_n210_n170#
+ m1_n1220_n5790# Vout Vout m1_n1220_n5790# m1_n1220_n5790# Vout Vout VSS m1_n210_n170#
+ sky130_fd_pr__nfet_01v8_GLZPWL
.ends

.subckt in_ring io_analog[10] vccd2 vssa2 vssd2 m2_1090872_693600# m3_601000_1115140#
+ m2_839106_693600# m2_633438_693600# m3_925294_1395900# m3_601000_944816# m2_798918_693600#
+ m2_609798_693600# m3_601000_1027514# m2_810738_693600# m3_1184520_714056# m2_1045956_693600#
+ m2_1151154_693600# m2_694902_693600# m3_1184520_1281890# m2_776460_693600# m2_953760_693600#
+ m2_1106238_693600# m2_1171248_693600# m2_631074_693600# m3_601000_1202766# m2_796554_693600#
+ m2_1002222_693600# m3_601000_1157180# m3_601000_1073100# m2_908844_693600# m2_973854_693600#
+ m2_1167702_693600# m2_1043592_693600# m3_601000_1069554# m3_1184520_1188922# analog_mux_0/SIG9
+ m2_651168_693600# m2_928938_693600# m2_1022316_693600# m2_993948_693600# m2_647622_693600#
+ m2_1063686_693600# m2_729180_693600# m2_930120_693600# m3_601000_705782# m3_1184520_708146#
+ m2_824922_693600# m2_794190_693600# m2_688992_693600# m2_906480_693600# m2_971490_693600#
+ m3_601000_1160726# m3_601000_728386# m3_1184520_1100078# m3_1184520_1057202# m2_667716_693600#
+ m3_601000_1200402# m3_1184520_1148046# m2_749274_693600# m2_950214_693600# m2_926574_693600#
+ m2_991584_693600# m3_1184520_717602# w_1135289_983102# m2_793008_693600# m2_769368_693600#
+ m2_970308_693600# m2_1040046_693600# a_1137371_982018# m2_946668_693600# m2_665352_693600#
+ m2_842652_693600# m2_1036500_693600# m3_601000_726022# m2_1077870_693600# m2_685446_693600#
+ m3_721194_1395900# m2_862746_693600# m2_1138152_693600# m2_1097964_693600# m2_923028_693600#
+ m2_787098_693600# m1_624380_1395640# m2_964398_693600# m2_1158246_693600# m3_601000_813648#
+ m2_683082_693600# m2_618072_693600# m3_1184520_1103624# m2_713814_693600# m2_860382_693600#
+ m2_1054230_693600# m3_601000_985474# m3_1184520_785172# m2_638166_693600# m2_733908_693600#
+ m2_1009314_693600# m3_1014394_1395900# m3_1184520_711692# m2_815466_693600# m2_1074324_693600#
+ m2_880476_693600# m2_699630_693600# m2_711450_693600# m2_876930_693600# m3_601000_699872#
+ m3_601000_771608# m2_1029408_693600# m2_1094418_693600# m2_937212_693600# m2_731544_693600#
+ m2_978582_693600# m3_601000_983110# m2_957306_693600# m2_751638_693600# m2_1027044_693600#
+ m2_833196_693600# m2_727998_693600# m2_998676_693600# m2_1092054_693600# m3_1183340_840430#
+ m3_1184520_705782# m3_1184520_741696# m2_829650_693600# m2_623982_693600# m2_894660_693600#
+ m2_1047138_693600# m2_602706_693600# m2_849744_693600# m2_1120422_693600# m2_1161792_693600#
+ m2_704358_693600# m2_975036_693600# m2_869838_693600# m2_806010_693600# m2_1140516_693600#
+ m2_871020_693600# m2_765822_693600# m2_1116876_693600# m2_1181886_693600# m2_847380_693600#
+ m3_601000_1117504# m2_1012860_693600# m2_620436_693600# m3_1184520_1013162# m2_891114_693600#
+ m2_826104_693600# m2_785916_693600# m2_867474_693600# m2_681900_693600# m2_1032954_693600#
+ m3_601000_702236# m2_722088_693600# m2_887568_693600# m3_601000_1159544# m2_718542_693600#
+ m2_989220_693600# m2_783552_693600# m3_601000_941270# m2_960852_693600# m2_1154700_693600#
+ m1_646350_1383430# m2_1030590_693600# m2_738636_693600# m2_1079052_693600# m2_915936_693600#
+ m2_980946_693600# m2_634620_693600# m2_1050684_693600# m3_1184520_699872# m2_811920_693600#
+ m2_675990_693600# m2_1099146_693600# m2_654714_693600# m2_1005768_693600# m2_1070778_693600#
+ m2_736272_693600# analog_mux_0/SEL0 m2_913572_693600# m2_1107420_693600# m2_1172430_693600#
+ m2_1148790_693600# m2_780006_693600# m2_674808_693600# m2_756366_693600# m2_933666_693600#
+ m3_601000_816012# m2_1127514_693600# m2_652350_693600# m2_1168884_693600# m3_601000_1199220#
+ m2_607434_693600# m2_1147608_693600# m2_878112_693600# m2_672444_693600# m2_1023498_693600#
+ m2_1019952_693600# m2_1125150_693600# m2_1084962_693600# m2_692538_693600# m2_627528_693600#
+ m2_910026_693600# m2_898206_693600# m2_774096_693600# m2_709086_693600# m2_804828_693600#
+ m2_668898_693600# analog_mux_0/SEL2 m2_605070_693600# m2_951396_693600# m2_1145244_693600#
+ m3_601000_696326# m2_700812_693600# m2_670080_693600# analog_mux_0/SIG11 m2_947850_693600#
+ m3_601000_987838# m3_1184520_787536# m2_1165338_693600# m5_930294_1395900# m2_690174_693600#
+ m2_625164_693600# a_606902_986681# m2_720906_693600# m3_1184520_1283072# m2_802464_693600#
+ m2_967944_693600# m2_1061322_693600# m3_1184520_744060# m2_1037682_693600# m3_774394_1395900#
+ m3_1184520_702236# m2_645258_693600# m2_1016406_693600# m2_822558_693600# m2_1081416_693600#
+ m2_1057776_693600# analog_mux_0/SIG3 m2_924210_693600# m2_788280_693600# analog_mux_0/GND
+ m2_965580_693600# m2_767004_693600# m2_1118058_693600# m2_1183068_693600# m2_944304_693600#
+ m2_1014042_693600# m2_820194_693600# m2_714996_693600# m2_985674_693600# m2_1179522_693600#
+ m2_610980_693600# m2_1034136_693600# m2_840288_693600# m2_659442_693600# m3_601000_940088#
+ m2_836742_693600# m2_1095600_693600# m5_766594_1395900# m3_601000_773972# m2_679536_693600#
+ m3_1184520_1280708# m2_962034_693600# m2_856836_693600# a_1137371_982518# m2_938394_693600#
+ analog_mux_0/SIG1 m2_752820_693600# m2_1103874_693600# m2_982128_693600# m3_601000_1028696#
+ m2_917118_693600# m2_958488_693600# m2_813102_693600# m2_677172_693600# m2_772914_693600#
+ m2_707904_693600# m2_1123968_693600# m2_854472_693600# m2_1048320_693600# m2_1089690_693600#
+ m2_697266_693600# m3_601000_1074282# m3_1184520_1193650# m2_809556_693600# m2_603888_693600#
+ m2_1068414_693600# m3_1184520_696326# m2_874566_693600# m3_601000_943634# m2_770550_693600#
+ m2_705540_693600# m3_601000_1026332# m2_1088508_693600# m2_1100328_693600# m2_725634_693600#
+ m2_996312_693600# m2_1141698_693600# m2_807192_693600# m2_790644_693600# m2_1066050_693600#
+ m2_902934_693600# m3_1184520_1058384# m3_601000_1201584# m2_745728_693600# m2_827286_693600#
+ m2_1086144_693600# m3_601000_1113958# m5_776894_1395900# m2_892296_693600# m2_641712_693600#
+ analog_mux_0/SIG0 m2_723270_693600# m2_888750_693600# m2_900570_693600# m2_661806_693600#
+ m2_949032_693600# m2_743364_693600# m2_920664_693600# m2_1114512_693600# m3_1184520_1056020#
+ m2_1155882_693600# m3_601000_1155998# m3_601000_1071918# m2_969126_693600# m2_763458_693600#
+ m3_1184520_716420# m2_940758_693600# analog_mux_0/SIG12 m2_1134606_693600# m2_865110_693600#
+ m2_759912_693600# m2_1010496_693600# m3_1183340_1234162# m2_1175976_693600# m3_826094_1395900#
+ m2_1006950_693600# m2_1071960_693600# m2_614526_693600# m2_885204_693600# m2_761094_693600#
+ m2_655896_693600# m2_1132242_693600# m3_1184524_1053656# m2_781188_693600# m2_716178_693600#
+ m4_930294_1395900# m2_612162_693600# m2_1152336_693600# m2_1128696_693600# m2_777642_693600#
+ m3_927794_1395900# m2_954942_693600# m2_1024680_693600# m3_1184520_1102442# m3_601000_812466#
+ m2_632256_693600# m2_797736_693600# m2_1003404_693600# m2_879294_693600# m3_601000_984292#
+ m2_628710_693600# m2_1044774_693600# m2_693720_693600# m5_818294_1395900# m2_858018_693600#
+ m2_899388_693600# m2_1105056_693600# m3_601000_709328# m2_754002_693600# m2_648804_693600#
+ m2_1064868_693600# m2_1170066_693600# m2_931302_693600# m3_601000_698690# m3_601000_770426#
+ m2_795372_693600# m2_1001040_693600# m3_1184520_1279526# m2_907662_693600# m2_701994_693600#
+ m2_972672_693600# m2_1166520_693600# m3_1184520_1192468# m2_927756_693600# m2_1021134_693600#
+ m2_992766_693600# m2_646440_693600# m5_919994_1395900# m2_823740_693600# m4_766594_1395900#
+ m2_1041228_693600# m2_666534_693600# m2_1017588_693600# m2_1082598_693600# m2_748092_693600#
+ m2_843834_693600# m2_925392_693600# m2_1119240_693600# m2_1184250_693600# m3_1184520_1190104#
+ m2_686628_693600# m2_904116_693600# m2_768186_693600# m2_863928_693600# m2_945486_693600#
+ m2_1139334_693600# m2_800100_693600# m2_664170_693600# m2_1110966_693600# m3_1111400_1392200#
+ m2_841470_693600# m2_1159428_693600# m2_684264_693600# m2_619254_693600# m5_828594_1395900#
+ m3_601000_1116322# m2_861564_693600# m2_1055412_693600# m2_1096782_693600# m3_1184520_715238#
+ m2_639348_693600# m2_816648_693600# m2_1075506_693600# m2_881658_693600# m2_1157064_693600#
+ m2_918300_693600# m2_712632_693600# m1_1149820_1377960# m2_983310_693600# m3_601000_701054#
+ m2_959670_693600# m1_1149820_1378460# m3_601000_1203948# m3_601000_1158362# m2_1177158_693600#
+ m4_776894_1395900# m2_732726_693600# m2_1008132_693600# m2_814284_693600# m2_979764_693600#
+ m2_1073142_693600# m3_601000_710510# m2_657078_693600# m3_601000_706964# m3_601000_817194#
+ m2_1028226_693600# m3_1184520_709328# m2_834378_693600# m2_999858_693600# m2_1093236_693600#
+ m3_1184520_698690# m2_936030_693600# m2_1069596_693600# m3_601000_729568# m2_730362_693600#
+ m3_1184520_1149228# m2_895842_693600# m2_1101510_693600# m2_1142880_693600# m2_956124_693600#
+ m2_750456_693600# m2_997494_693600# m2_1121604_693600# m2_746910_693600# m2_1162974_693600#
+ m3_601000_704600# m2_976218_693600# m2_601524_693600# m3_601000_727204# m2_872202_693600#
+ m2_642894_693600# m2_848562_693600# m2_621618_693600# m2_703176_693600# m3_930294_1395900#
+ m2_662988_693600# m2_868656_693600# m2_764640_693600# m2_1115694_693600# m3_1184520_1104806#
+ m3_601000_769244# m2_941940_693600# m3_601000_695144# m3_771894_1395900# m2_719724_693600#
+ m2_1135788_693600# m3_601000_986656# m2_784734_693600# m3_1184520_786354# m2_866292_693600#
+ m3_1184520_712874# m2_1031772_693600# m4_818294_1395900# m2_845016_693600# m2_739818_693600#
+ m2_886386_693600# m2_741000_693600# m2_635802_693600# m2_1051866_693600# m3_1184520_701054#
+ m2_717360_693600# m3_1066100_1382200# m2_782370_693600# m2_1112148_693600# m2_737454_693600#
+ m3_1184520_710510# m2_914754_693600# m2_1108602_693600# m2_1173612_693600# analog_mux_0/SIG2
+ m4_919994_1395900# m2_1149972_693600# m3_766594_1395900# m3_1184520_706964# m3_601000_730750#
+ m3_1184520_742878# m2_757548_693600# m2_934848_693600# m2_859200_693600# m2_653532_693600#
+ m2_1004586_693600# m2_735090_693600# m2_629892_693600# m2_830832_693600# m2_912390_693600#
+ m2_608616_693600# m2_673626_693600# m2_755184_693600# m2_649986_693600# m2_850926_693600#
+ m2_932484_693600# m3_601000_772790# m2_1126332_693600# m3_1184520_704600# m3_1184520_740514#
+ m3_1183340_1244162# m2_911208_693600# m2_775278_693600# m4_828594_1395900# m3_601000_1031060#
+ m2_606252_693600# m2_952578_693600# m2_1146426_693600# m2_671262_693600# m2_1042410_693600#
+ m2_1018770_693600# m2_1083780_693600# m3_1174000_874700# m2_897024_693600# m2_691356_693600#
+ m2_626346_693600# m2_803646_693600# m2_1062504_693600# m2_1038864_693600# m2_1144062_693600#
+ m3_601000_703418# m2_687810_693600# a_606902_945081# m3_1184520_695144# m3_776894_1395900#
+ m3_601000_942452# m2_905298_693600# m2_1058958_693600# m2_1164156_693600# m2_789462_693600#
+ m2_990402_693600# m2_801282_693600# m2_966762_693600# m2_1060140_693600# m2_644076_693600#
+ m2_1015224_693600# m2_821376_693600# m2_986856_693600# m2_1080234_693600# m2_1056594_693600#
+ m2_817830_693600# m2_882840_693600# m3_601000_1112776# m2_1035318_693600# m3_1183340_830430#
+ m2_1076688_693600# m2_943122_693600# m2_837924_693600# m2_919482_693600# m2_984492_693600#
+ m2_1178340_693600# m2_963216_693600# m3_823594_1395900# m2_939576_693600# m2_658260_693600#
+ m3_601000_1070736# m2_835560_693600# m2_1053048_693600# m2_678354_693600# m2_855654_693600#
+ m2_1049502_693600# m2_1102692_693600# m3_601000_697508# m2_698448_693600# m2_710268_693600#
+ m3_1184520_1054838# m2_875748_693600# m3_1184520_788718# m2_771732_693600# m2_706722_693600#
+ m2_977400_693600# m2_1122786_693600# m2_853290_693600# m3_818294_1395900# m2_696084_693600#
+ m2_832014_693600# m2_726816_693600# m2_808374_693600# m2_791826_693600# m2_1067232_693600#
+ m3_1184520_1101260# m3_1184520_703418# m2_873384_693600# m2_622800_693600# m2_852108_693600#
+ m2_828468_693600# m2_1087326_693600# m2_893478_693600# m2_724452_693600# m2_995130_693600#
+ analog_mux_0/SEL1 m2_889932_693600# m3_919994_1395900# m3_601000_708146# m2_901752_693600#
+ m2_1160610_693600# m2_1136970_693600# m3_1184520_1278344# analog_mux_0/SIG4 m2_744546_693600#
+ m3_1184520_1191286# m2_921846_693600# m2_1180704_693600# analog_mux_0/OUT m2_640530_693600#
+ m2_616890_693600# m2_846198_693600# m2_660624_693600# m2_1011678_693600# m2_742182_693600#
+ m2_636984_693600# m3_601000_814830# m2_1113330_693600# m3_1148600_1374300# m2_615708_693600#
+ analog_mux_0/SEL3 vdda2 m2_680718_693600# m2_762276_693600# m3_828594_1395900# m2_1133424_693600#
+ m3_601000_1029878# m2_758730_693600# m2_1109784_693600# m2_1174794_693600# m2_988038_693600#
+ m2_613344_693600# m2_1153518_693600# m2_884022_693600# m2_819012_693600# m2_1129878_693600#
+ m2_778824_693600# m2_1025862_693600# m2_1131060_693600# m3_1184520_697508#
Xdiode_connected_nmos_6 m3_1148600_1374300# m1_1149820_1377960# analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_7 m1_1149820_1377960# analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
Xanalog_mux_0 analog_mux_0/OUT vdda2 analog_mux_0/SIG0 analog_mux_0/SIG1 analog_mux_0/SIG2
+ analog_mux_0/SIG3 analog_mux_0/SIG4 analog_mux_0/SIG5 analog_mux_0/SIG6 analog_mux_0/SIG7
+ vdda2 analog_mux_0/SIG9 analog_mux_0/GND analog_mux_0/SIG11 analog_mux_0/SIG12 analog_mux_0/SIG13
+ analog_mux_0/SIG14 analog_mux_0/SIG15 analog_mux_0/SEL0 analog_mux_0/SEL1 analog_mux_0/SEL2
+ analog_mux_0/SEL3 analog_mux_0/GND analog_mux
XOTA_fingers_031123_NON_FLAT_0 io_analog[10] m1_624380_1395640# vccd2 constant_gm_fingers_0/Vout
+ m1_646350_1383430# analog_mux_0/GND OTA_fingers_031123_NON_FLAT
Xdiode_connected_nmos_0 vccd2 m1_624380_1395640# analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_1 m1_624380_1395640# analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_2 m1_646350_1383430# analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_4 m1_1149820_1378460# analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
XOTA_MULT_GM_0 m3_1148600_1374300# m1_1149820_1377960# m1_1149820_1378460# m3_1148600_1374300#
+ m3_1066100_1382200# analog_mux_0/GND OTA_MULT_GM
Xdiode_connected_nmos_3 vccd2 m1_646350_1383430# analog_mux_0/GND diode_connected_nmos
Xconstant_gm_fingers_0 constant_gm_fingers_0/Vout vccd2 analog_mux_0/GND constant_gm_fingers
Xdiode_connected_nmos_5 m3_1148600_1374300# m1_1149820_1378460# analog_mux_0/GND diode_connected_nmos
X0 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=7.44e+13p ps=5.2976e+08u w=5e+06u l=500000u
X1 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X2 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=1.3679e+14p pd=1.00302e+09u as=1.595e+13p ps=1.1638e+08u w=5e+06u l=500000u
X3 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X4 w_1135289_983102# a_1137371_982018# a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=3.81686e+14p pd=3.65032e+09u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X5 w_1135289_983102# a_1137371_982518# a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X6 analog_mux_0/SIG7 a_612871_959293# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X7 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X8 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=4.54e+13p pd=3.1816e+08u as=0p ps=0u w=5e+06u l=500000u
X9 a_1137916_978034# a_1137916_978034# analog_mux_0/SIG13 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=1.105e+13p ps=7.674e+07u w=2.5e+06u l=500000u
X10 w_1135289_983102# a_1137916_978034# a_1137916_978034# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X11 analog_mux_0/SIG14 a_1137371_982518# a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.83e+13p pd=1.2732e+08u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=500000u
X12 analog_mux_0/GND analog_mux_0/SIG6 a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=7.17928e+14p pd=5.06904e+09u as=2.32e+13p ps=1.6928e+08u w=5e+06u l=1e+06u
X13 a_615374_964626# a_606902_945081# a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=5.8e+12p pd=4.232e+07u as=0p ps=0u w=5e+06u l=500000u
X14 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_618579_965827# a_606902_986681# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.395e+13p ps=9.558e+07u w=5e+06u l=500000u
X16 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=3.235e+13p pd=2.2294e+08u as=0p ps=0u w=5e+06u l=500000u
X17 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_618579_965827# a_606902_945081# a_615374_964626# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.685e+13p ps=3.2874e+08u w=5e+06u l=500000u
X21 vdda2 a_606902_945081# a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=3.18606e+14p pd=2.87548e+09u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X22 analog_mux_0/SIG5 a_612871_959293# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X23 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X24 a_1137371_982518# a_1137371_982518# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X25 a_1137371_982518# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X26 analog_mux_0/GND analog_mux_0/GND a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X27 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X28 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X29 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X30 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X31 analog_mux_0/SIG14 a_1131722_982955# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X32 a_1137371_982018# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X33 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X34 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X35 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X36 vdda2 a_625084_965506# analog_mux_0/SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.075e+13p ps=1.383e+08u w=5e+06u l=1e+06u
X37 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X38 analog_mux_0/GND analog_mux_0/GND a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X39 a_618579_965827# a_606902_986681# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X40 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X41 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X42 analog_mux_0/GND analog_mux_0/GND a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X43 w_1135289_983102# a_1137916_978034# a_1137916_978034# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X44 a_1137459_979540# a_1137371_982018# a_1137271_985458# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X45 a_606902_945081# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X46 analog_mux_0/GND analog_mux_0/GND a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X47 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.83e+13p pd=1.2732e+08u as=0p ps=0u w=5e+06u l=1e+06u
X48 a_1137371_982018# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X49 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X50 a_606902_986681# a_606902_986681# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X51 analog_mux_0/SIG5 a_606902_986681# a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X52 a_615374_964626# a_606902_945081# a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X53 a_606902_986681# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X54 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X55 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X56 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=2.555e+13p pd=1.8022e+08u as=0p ps=0u w=5e+06u l=1e+06u
X57 analog_mux_0/GND analog_mux_0/GND a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X58 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X59 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X60 analog_mux_0/GND analog_mux_0/GND a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X61 a_618579_965827# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X62 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X63 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X64 a_618579_965827# a_606902_945081# a_615374_964626# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X65 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X66 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X67 analog_mux_0/SIG14 a_1137371_982518# a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X68 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X69 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X70 a_1137371_982518# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X71 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.6e+12p ps=6.5e+07u w=1.25e+06u l=1e+06u
X72 a_1137459_979540# a_1137371_982018# a_1137271_985458# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X73 a_606902_986681# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X74 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X75 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X76 analog_mux_0/GND analog_mux_0/GND a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X77 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X78 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X79 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X80 a_618579_965827# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X81 analog_mux_0/GND a_1138059_976036# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X82 a_630040_965691# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X83 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X84 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X85 vdda2 a_606902_986681# a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X86 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X87 vdda2 a_625084_965506# a_625084_965506# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X88 a_618579_965827# a_606902_986681# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X89 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X90 a_606902_986681# a_606902_986681# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X91 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X92 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X93 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X94 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X95 analog_mux_0/SIG15 a_1131722_982955# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X96 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X97 vdda2 a_606902_986681# a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X98 w_1135289_983102# a_1137916_978034# analog_mux_0/SIG13 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.51e+13p ps=1.7004e+08u w=5e+06u l=1e+06u
X99 analog_mux_0/SIG5 a_606902_986681# a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X100 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X101 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X102 analog_mux_0/GND a_1138059_976036# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X103 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X104 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X105 a_606902_986681# a_606902_986681# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X106 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X107 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X108 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X109 w_1135289_983102# a_1137916_978034# analog_mux_0/SIG13 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X110 a_1137459_979540# a_1137371_982018# a_1137271_985458# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X111 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X112 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X113 analog_mux_0/SIG6 a_625084_965506# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X114 w_1135289_983102# a_1137916_978034# a_1137916_978034# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X115 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X116 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X117 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X118 analog_mux_0/GND a_1138059_976036# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X119 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X120 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X121 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X122 a_1137916_978034# analog_mux_0/SIG13 a_1138059_976036# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X123 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X124 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X125 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X126 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X127 a_1137916_978034# analog_mux_0/SIG13 a_1138059_976036# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X128 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X129 analog_mux_0/SIG15 a_1131722_982955# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X130 analog_mux_0/SIG7 a_612871_959293# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X131 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X132 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X133 analog_mux_0/GND analog_mux_0/GND a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X134 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X135 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X136 vdda2 a_625084_965506# analog_mux_0/SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X137 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X138 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X139 analog_mux_0/GND analog_mux_0/SIG6 a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X140 a_630040_965691# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X141 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X142 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X143 a_1137371_982018# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X144 a_606902_945081# a_606902_945081# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X145 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X146 a_630040_965691# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X147 analog_mux_0/GND analog_mux_0/GND a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X148 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X149 a_1131722_982955# analog_mux_0/SIG14 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X150 w_1135289_983102# a_1137916_978034# a_1137916_978034# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X151 vdda2 a_606902_945081# a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X152 analog_mux_0/GND analog_mux_0/SIG6 a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X153 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X154 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X155 a_625084_965506# analog_mux_0/SIG6 a_630040_965691# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=7.25e+12p pd=5.348e+07u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X156 analog_mux_0/GND analog_mux_0/GND a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X157 a_606902_945081# a_606902_945081# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X158 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X159 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X160 analog_mux_0/SIG15 a_1131722_982955# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X161 a_625084_965506# a_625084_965506# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X162 a_625084_965506# analog_mux_0/SIG6 a_630040_965691# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X163 vdda2 a_606902_945081# a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X164 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X165 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X166 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X167 a_606902_945081# a_606902_945081# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X168 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X169 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X170 analog_mux_0/GND analog_mux_0/GND a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X171 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X172 a_618579_965827# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X173 a_606902_945081# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X174 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X175 a_1137371_982018# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X176 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X177 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X178 a_606902_986681# a_606902_986681# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X179 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X180 a_606902_986681# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X181 analog_mux_0/GND analog_mux_0/GND a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X182 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X183 vdda2 a_625084_965506# a_625084_965506# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X185 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X186 vdda2 a_606902_986681# a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X187 a_1137916_978034# analog_mux_0/SIG13 a_1138059_976036# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X188 analog_mux_0/GND analog_mux_0/GND a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X189 a_606902_945081# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X190 analog_mux_0/SIG15 a_1131722_982955# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X191 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X192 a_606902_986681# a_606902_986681# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X193 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X194 analog_mux_0/GND analog_mux_0/GND a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X195 a_606902_986681# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X196 a_630040_965691# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X197 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X198 vdda2 a_606902_986681# a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X199 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X200 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X201 a_612871_959293# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X202 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X203 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X204 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X205 analog_mux_0/SIG6 a_625084_965506# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X206 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X207 analog_mux_0/SIG14 a_1137371_982518# a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X208 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X209 a_618579_965827# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X210 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X211 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 w_1135289_983102# a_1137371_982518# a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X213 a_630040_965691# analog_mux_0/SIG6 a_625084_965506# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X214 w_1135289_983102# a_1137371_982518# a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X215 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
R0 vssa2 analog_mux_0/GND sky130_fd_pr__res_generic_m3 w=7.45e+07u l=2.6e+06u
X216 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X217 a_1137371_982518# a_1137371_982518# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X218 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X219 analog_mux_0/SIG7 a_612871_959293# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X220 a_1137916_978034# a_1137916_978034# analog_mux_0/SIG13 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X221 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X222 a_606902_945081# a_606902_945081# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X223 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X224 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X225 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X226 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X227 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X228 a_625084_965506# a_625084_965506# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X229 analog_mux_0/GND analog_mux_0/SIG6 a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X230 a_1137459_979540# a_1137371_982018# a_1137271_985458# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X231 analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X232 a_612871_959293# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X233 analog_mux_0/GND a_1138059_976036# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X234 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X235 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X236 w_1135289_983102# a_1137371_982518# a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X237 analog_mux_0/GND analog_mux_0/GND a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X238 w_1135289_983102# a_1137371_982018# a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X239 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X240 analog_mux_0/GND analog_mux_0/GND a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X241 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
R1 analog_mux_0/GND m3_1174000_874700# sky130_fd_pr__res_generic_m3 w=7.7e+07u l=5e+06u
X242 vdda2 a_606902_945081# a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X243 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X244 a_1137371_982518# a_1137371_982518# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X245 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X246 a_606902_945081# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X247 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X248 a_1137371_982518# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X249 vdda2 a_625084_965506# analog_mux_0/SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X250 a_606902_945081# a_606902_945081# vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X251 analog_mux_0/SIG14 a_1137371_982518# a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X252 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X253 w_1135289_983102# a_1137916_978034# analog_mux_0/SIG13 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X254 analog_mux_0/GND analog_mux_0/GND a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X255 a_1137459_979540# a_1137371_982018# a_1137271_985458# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X256 vdda2 a_606902_945081# a_606902_945081# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X257 a_606902_945081# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X258 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X259 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X260 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X261 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X262 analog_mux_0/SIG14 a_1137371_982518# a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X263 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X264 analog_mux_0/GND analog_mux_0/GND a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X265 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X266 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X267 a_1137371_982518# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X268 a_618579_965827# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X269 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X270 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X271 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X272 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X273 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X274 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X275 w_1135289_983102# a_1137916_978034# analog_mux_0/SIG13 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X276 a_618579_965827# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X277 vdda2 a_625084_965506# a_625084_965506# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X278 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
R2 analog_mux_0/GND m3_1111400_1392200# sky130_fd_pr__res_generic_m4 w=2.75e+07u l=2.8e+06u
X279 w_1135289_983102# a_1137916_978034# a_1137916_978034# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X280 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X281 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X282 a_1137371_982518# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X283 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X284 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X285 w_1135289_983102# a_1137916_978034# a_1137916_978034# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X286 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X287 analog_mux_0/SIG14 a_1137371_982518# a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X288 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X289 analog_mux_0/GND analog_mux_0/GND a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X290 a_1137459_979540# a_1137371_982018# a_1137271_985458# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X291 a_1131722_982955# analog_mux_0/SIG14 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X292 analog_mux_0/SIG14 a_1131722_982955# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X293 analog_mux_0/SIG6 a_625084_965506# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X294 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X295 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X296 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X297 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X298 a_1137916_978034# analog_mux_0/SIG13 a_1138059_976036# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X299 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X300 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X301 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X302 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X303 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X304 a_1137371_982018# a_1137371_982018# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X305 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X306 analog_mux_0/GND analog_mux_0/GND a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X307 analog_mux_0/SIG7 a_612871_959293# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X308 w_1135289_983102# a_1137371_982018# a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X309 a_1137371_982018# a_1137371_982018# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X310 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X311 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X312 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X313 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X314 analog_mux_0/GND analog_mux_0/SIG6 a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X315 analog_mux_0/GND analog_mux_0/SIG6 a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X316 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X317 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X318 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X319 w_1135289_983102# a_1137916_978034# analog_mux_0/SIG13 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X320 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X321 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X322 a_625084_965506# a_625084_965506# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X323 analog_mux_0/GND analog_mux_0/SIG6 a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X324 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X325 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X326 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X327 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X328 w_1135289_983102# a_1137371_982018# a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X329 vdda2 a_615374_964626# a_615374_964626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X330 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X331 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X332 analog_mux_0/SIG6 a_625084_965506# a_625084_965506# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X333 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X334 a_1137371_982018# a_1137371_982018# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X335 a_625084_965506# analog_mux_0/SIG6 a_630040_965691# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X336 a_1137371_982018# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X337 a_1137916_978034# analog_mux_0/SIG13 a_1138059_976036# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X338 w_1135289_983102# a_1137916_978034# analog_mux_0/SIG13 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X339 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X340 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X341 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X342 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X343 a_618579_965827# a_606902_945081# a_615374_964626# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X344 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X345 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X346 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X347 a_606902_986681# analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X348 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X349 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X350 a_1137916_978034# analog_mux_0/SIG13 a_1138059_976036# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X351 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X352 a_618579_965827# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X353 w_1135289_983102# a_1137271_985458# a_1137271_985458# w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X354 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X355 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X356 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X357 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X358 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X359 a_1137371_982518# a_1137371_982518# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X360 analog_mux_0/SIG5 a_606902_986681# a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X361 a_615374_964626# a_606902_945081# a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
R3 vssd2 analog_mux_0/GND sky130_fd_pr__res_generic_m3 w=7.55e+07u l=1e+07u
X362 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X363 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X364 vdda2 a_606902_986681# a_606902_986681# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X365 analog_mux_0/SIG5 a_612871_959293# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X366 w_1135289_983102# a_1137371_982518# a_1137371_982518# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X367 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X368 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X369 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X370 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X371 a_615374_964626# a_606902_945081# a_618579_965827# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X372 vdda2 a_615374_964626# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X373 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X374 w_1135289_983102# a_1137271_985458# analog_mux_0/SIG14 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X375 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X376 a_1137371_982018# a_1137371_982018# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X377 analog_mux_0/SIG14 a_1137371_982518# a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X378 a_630040_965691# analog_mux_0/SIG6 a_625084_965506# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X379 analog_mux_0/SIG5 a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X380 a_630040_965691# analog_mux_0/SIG6 a_625084_965506# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X381 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X382 a_1137459_979540# a_1137371_982018# a_1137271_985458# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X383 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X384 analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X385 a_615374_964626# a_615374_964626# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X386 w_1135289_983102# a_1137371_982018# a_1137371_982018# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X387 analog_mux_0/GND analog_mux_0/SIG13 a_1137459_979540# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X388 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X389 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X390 a_1137371_982518# a_1137371_982518# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X391 a_618579_965827# a_606902_986681# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X392 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X393 w_1135289_983102# analog_mux_0/SIG14 analog_mux_0/SIG15 w_1135289_983102# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X394 a_625084_965506# a_625084_965506# analog_mux_0/SIG6 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X395 a_1137371_982018# a_1137371_982018# w_1135289_983102# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
.ends

.subckt lvs gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12] gpio_analog[13]
+ gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[17] gpio_analog[1] gpio_analog[2]
+ gpio_analog[3] gpio_analog[4] gpio_analog[5] gpio_analog[6] gpio_analog[7] gpio_analog[8]
+ gpio_analog[9] gpio_noesd[0] gpio_noesd[10] gpio_noesd[11] gpio_noesd[12] gpio_noesd[13]
+ gpio_noesd[14] gpio_noesd[15] gpio_noesd[16] gpio_noesd[17] gpio_noesd[1] gpio_noesd[2]
+ gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6] gpio_noesd[7] gpio_noesd[8]
+ gpio_noesd[9] io_analog[0] io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5]
+ io_analog[6] io_analog[7] io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1]
+ io_clamp_high[2] io_clamp_low[0] io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10]
+ io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26]
+ io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0]
+ io_in_3v3[10] io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[14] io_in_3v3[15]
+ io_in_3v3[16] io_in_3v3[17] io_in_3v3[18] io_in_3v3[19] io_in_3v3[1] io_in_3v3[20]
+ io_in_3v3[21] io_in_3v3[22] io_in_3v3[23] io_in_3v3[24] io_in_3v3[25] io_in_3v3[26]
+ io_in_3v3[2] io_in_3v3[3] io_in_3v3[4] io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8]
+ io_in_3v3[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2
+ user_irq[0] user_irq[1] user_irq[2] vccd1 vdda1 vssa1 vssd1 wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xin_ring_0 in_ring_0/io_analog[10] in_ring_0/vccd2 in_ring_0/vssa2 in_ring_0/vssd2
+ la_oenb[102] io_in[16] la_oenb[31] wbs_dat_o[5] io_clamp_low[0] gpio_noesd[13] la_data_out[20]
+ wbs_dat_i[0] io_out[18] la_oenb[23] io_in_3v3[4] la_data_in[90] la_oenb[119] wbs_adr_i[23]
+ io_out[13] la_data_in[14] la_data_in[64] la_data_in[107] la_data_out[125] wbs_adr_i[5]
+ io_in_3v3[14] la_oenb[19] la_oenb[77] io_out[15] io_in_3v3[17] la_data_out[51] la_oenb[69]
+ la_data_out[124] la_data_out[89] io_oeb[17] gpio_noesd[5] gpio_analog[14] wbs_dat_o[10]
+ la_data_in[57] la_data_out[83] la_data_out[75] wbs_dat_o[9] la_data_in[95] la_oenb[0]
+ la_data_out[57] io_out[24] io_oeb[2] la_oenb[27] la_data_in[19] wbs_dat_i[21] la_oenb[50]
+ la_data_in[69] gpio_noesd[8] io_in[23] gpio_noesd[3] io_out[9] wbs_dat_i[15] io_out[14]
+ io_out[11] la_data_out[6] la_data_in[63] la_data_out[56] la_oenb[74] io_oeb[4] vdda1
+ la_oenb[18] la_data_in[12] la_oenb[68] la_data_out[88] gpio_analog[0] la_data_in[62]
+ wbs_dat_o[14] la_oenb[32] la_data_out[87] io_oeb[23] la_data_in[99] wbs_dat_i[20]
+ io_analog[7] la_data_out[38] la_data_in[116] la_oenb[104] la_data_out[55] la_data_in[17]
+ io_analog[9] la_data_in[67] la_oenb[121] io_out[21] wbs_dat_o[19] wbs_adr_i[2] io_out[10]
+ wbs_dat_i[28] la_oenb[37] la_data_out[92] io_in[19] io_in_3v3[6] wbs_adr_i[7] la_data_in[2]
+ la_oenb[79] io_analog[3] io_out[3] la_data_in[25] la_data_in[98] la_data_out[43]
+ wbs_dat_i[24] wbs_dat_o[27] la_data_out[42] io_oeb[25] io_in[22] la_data_out[85]
+ la_oenb[103] la_data_out[59] la_data_out[1] la_data_in[71] io_oeb[19] la_data_in[65]
+ la_data_in[7] la_oenb[84] la_data_in[30] la_data_out[0] la_oenb[76] la_data_in[103]
+ vssa1 io_in[2] io_in[5] la_data_in[29] wbs_dat_i[3] la_data_out[47] la_data_out[90]
+ wb_rst_i la_oenb[34] la_data_in[111] la_oenb[122] wbs_dat_o[25] la_data_in[70] la_data_out[40]
+ la_data_out[22] la_oenb[116] la_oenb[40] la_data_in[11] la_data_in[110] user_irq[0]
+ la_data_in[34] gpio_noesd[9] la_oenb[80] wbs_dat_o[2] io_oeb[8] la_data_out[46]
+ la_data_in[28] la_oenb[16] la_oenb[39] wbs_dat_i[19] la_data_out[86] io_in[25] wbs_dat_o[30]
+ la_data_out[45] io_in_3v3[15] wbs_dat_o[29] la_data_in[74] la_data_in[16] io_out[20]
+ la_data_in[66] la_oenb[120] io_analog[8] la_oenb[85] la_data_out[3] la_data_out[99]
+ la_data_out[53] la_oenb[71] wbs_adr_i[6] la_data_out[91] io_in_3v3[1] la_data_in[24]
+ wbs_dat_o[17] la_data_in[105] wbs_dat_o[11] la_oenb[78] la_data_in[97] la_oenb[2]
+ gpio_analog[6] la_oenb[52] la_data_out[107] la_oenb[125] la_data_in[119] la_data_in[15]
+ wbs_dat_i[17] la_data_out[8] la_data_out[58] io_in_3v3[21] la_data_in[113] wbs_adr_i[11]
+ la_oenb[124] io_oeb[14] wbs_we_i la_oenb[118] la_oenb[42] wbs_dat_o[16] la_oenb[83]
+ la_oenb[82] la_data_out[112] la_data_in[101] wbs_dat_i[22] wbs_adr_i[4] la_oenb[51]
+ la_data_out[48] la_data_out[13] wbs_adr_i[27] la_data_in[22] wbs_dat_o[15] gpio_analog[4]
+ wbs_cyc_i la_data_out[63] la_data_in[118] io_out[26] wbs_dat_o[24] wbs_adr_i[16]
+ gpio_analog[15] la_data_out[62] gpio_noesd[12] io_out[6] la_oenb[123] io_analog[4]
+ wbs_dat_o[21] wbs_dat_o[3] gpio_analog[12] wbs_dat_i[30] io_oeb[13] la_data_out[21]
+ la_data_in[68] la_data_out[94] io_oeb[5] la_oenb[87] io_clamp_high[2] io_out[1]
+ wbs_adr_i[9] la_oenb[81] la_data_in[27] la_data_in[100] la_data_out[93] gpio_analog[10]
+ la_oenb[55] la_data_out[17] VSUBS la_data_out[67] la_data_out[11] la_data_out[110]
+ user_irq[1] la_data_out[61] la_data_in[81] la_data_out[26] wbs_dat_o[28] la_data_in[73]
+ la_oenb[127] wbs_dat_o[0] la_oenb[86] la_data_in[32] wbs_adr_i[13] io_oeb[20] la_data_in[31]
+ la_data_in[104] io_analog[6] gpio_noesd[15] wbs_dat_o[18] io_in[13] la_data_out[66]
+ la_oenb[36] gpio_analog[1] la_oenb[59] gpio_analog[8] la_data_out[7] la_data_out[106]
+ la_data_in[72] io_in[18] la_oenb[53] la_data_out[65] la_data_out[24] wbs_adr_i[18]
+ la_data_in[13] wbs_dat_o[26] la_data_in[112] la_data_in[36] la_oenb[90] la_data_out[102]
+ wbs_dat_o[23] gpio_noesd[10] io_oeb[12] la_data_out[23] wbs_ack_o la_data_out[96]
+ io_in[0] la_oenb[41] io_in_3v3[20] la_data_out[12] wbs_adr_i[26] io_oeb[18] la_data_in[102]
+ la_data_out[105] wbs_dat_o[31] la_data_in[76] la_data_in[117] la_oenb[22] la_data_in[18]
+ la_oenb[95] la_oenb[49] io_oeb[9] io_in[14] la_data_out[5] la_data_out[28] la_data_out[101]
+ io_out[16] io_analog[6] la_oenb[46] wbs_adr_i[8] gpio_analog[7] wbs_adr_i[31] la_oenb[45]
+ la_data_in[49] wbs_dat_o[13] la_oenb[62] la_oenb[4] la_oenb[54] la_data_out[109]
+ io_in[9] la_data_in[121] io_oeb[15] io_in[17] la_data_out[68] la_data_out[10] io_out[4]
+ la_data_out[60] gpio_analog[16] la_data_in[115] la_data_in[39] la_data_out[9] la_data_in[80]
+ vdda1 la_oenb[126] io_clamp_high[1] la_data_in[79] la_data_out[97] wbs_dat_i[1]
+ la_oenb[44] la_oenb[9] wbs_adr_i[12] la_data_out[114] gpio_noesd[2] la_data_out[15]
+ wbs_adr_i[29] io_analog[4] wbs_sel_i[0] la_data_in[120] la_data_out[113] la_data_out[14]
+ io_clamp_high[0] la_data_out[64] la_data_in[84] io_in[10] io_oeb[21] wbs_dat_i[5]
+ la_data_in[20] la_data_in[78] la_data_in[43] io_out[19] wbs_dat_i[4] la_oenb[89]
+ wbs_dat_o[22] io_analog[5] la_data_in[37] la_oenb[48] la_oenb[106] gpio_noesd[17]
+ la_oenb[7] wbs_adr_i[10] la_data_out[95] la_data_in[125] la_oenb[57] io_in_3v3[26]
+ io_out[22] la_data_out[19] la_data_out[77] io_in_3v3[13] la_data_in[51] wbs_adr_i[25]
+ la_data_out[69] la_data_in[124] io_out[12] la_oenb[56] la_data_in[83] la_data_in[75]
+ wbs_dat_i[9] io_analog[4] la_data_out[27] io_analog[6] la_oenb[88] wbs_adr_i[15]
+ la_data_in[82] la_data_out[100] la_data_in[6] la_data_in[33] la_data_in[56] la_oenb[110]
+ user_irq[2] io_in_3v3[12] wbs_dat_o[20] la_data_in[50] la_oenb[11] la_oenb[38] la_oenb[61]
+ la_data_out[116] la_oenb[20] wbs_dat_i[14] la_data_out[108] vssa1 la_data_out[32]
+ la_data_in[122] wbs_adr_i[20] wbs_dat_i[2] io_analog[5] io_in_3v3[16] la_data_in[38]
+ la_oenb[92] la_data_out[104] io_in[4] wbs_dat_i[7] la_data_out[25] la_data_out[98]
+ la_oenb[43] la_data_out[121] la_data_in[54] wbs_adr_i[28] io_analog[0] la_data_out[72]
+ io_out[25] la_oenb[65] io_analog[1] gpio_noesd[7] io_in[15] la_data_in[127] io_analog[6]
+ la_oenb[1] la_data_out[79] la_oenb[24] la_data_out[71] la_oenb[97] gpio_analog[17]
+ wbs_dat_i[12] io_in[24] gpio_noesd[14] la_data_in[85] io_in_3v3[3] la_data_out[30]
+ la_data_in[77] la_data_out[103] io_oeb[0] la_data_in[59] la_oenb[96] io_in_3v3[23]
+ la_data_in[1] io_oeb[11] la_oenb[47] la_oenb[105] la_data_out[117] la_oenb[64] la_oenb[6]
+ la_data_out[76] la_data_out[111] la_oenb[5] la_data_in[123] io_oeb[24] la_data_out[70]
+ wb_clk_i io_out[23] la_data_in[41] wbs_dat_i[8] la_data_out[34] wbs_sel_i[2] wbs_dat_i[25]
+ io_analog[4] wbs_adr_i[14] la_data_in[40] la_oenb[10] la_oenb[109] io_oeb[10] io_oeb[22]
+ la_oenb[60] io_oeb[26] io_clamp_low[2] wbs_adr_i[30] la_data_out[115] io_in_3v3[19]
+ la_data_out[16] io_in[6] la_data_out[39] io_oeb[3] la_data_in[86] io_analog[5] la_data_out[33]
+ la_oenb[3] la_data_in[45] la_data_in[4] wbs_dat_i[6] la_oenb[91] io_in[1] wbs_dat_i[29]
+ io_analog[2] la_oenb[15] la_oenb[108] la_data_in[3] io_in[3] la_data_in[53] la_oenb[107]
+ la_data_in[126] gpio_analog[9] io_analog[4] la_data_out[119] io_analog[6] io_out[2]
+ gpio_noesd[16] io_out[5] la_oenb[8] la_oenb[58] la_data_out[37] wbs_dat_i[11] la_data_out[78]
+ la_data_out[2] wbs_dat_o[4] la_data_out[29] la_data_out[52] wbs_adr_i[0] wbs_adr_i[17]
+ la_data_in[8] wbs_dat_i[10] la_data_in[35] la_data_in[58] io_in_3v3[22] la_oenb[112]
+ io_in_3v3[2] io_in_3v3[5] vdda1 la_data_in[52] la_oenb[13] io_analog[5] gpio_noesd[11]
+ wbs_stb_i la_oenb[63] la_data_out[118] wbs_dat_i[16] la_data_in[89] la_data_out[82]
+ la_oenb[100] vssd1 la_data_in[48] wbs_adr_i[22] wbs_sel_i[3] la_oenb[21] la_oenb[94]
+ la_data_in[88] la_oenb[117] io_in_3v3[25] wbs_adr_i[21] gpio_analog[13] io_in_3v3[0]
+ io_analog[6] io_in[20] la_data_out[50] la_oenb[93] la_data_out[123] la_oenb[17]
+ la_data_out[74] la_data_in[21] la_oenb[67] la_data_in[94] wbs_dat_o[8] la_data_out[81]
+ la_oenb[26] la_data_out[73] la_oenb[99] la_data_in[93] la_oenb[25] la_data_in[44]
+ io_oeb[16] la_data_in[87] vssa1 la_oenb[98] la_data_in[61] la_data_out[31] la_data_out[54]
+ la_oenb[72] la_data_out[127] la_oenb[66] io_clamp_low[1] la_data_in[60] wbs_dat_o[12]
+ io_out[17] la_oenb[30] la_data_in[92] wbs_dat_i[18] la_data_out[36] la_data_in[91]
+ la_data_in[106] io_in[26] wbs_adr_i[24] wbs_dat_i[27] io_in_3v3[9] la_data_in[42]
+ io_oeb[6] la_oenb[12] wbs_dat_i[26] la_oenb[70] la_oenb[111] la_oenb[35] io_analog[5]
+ wbs_dat_i[23] la_oenb[29] la_data_in[0] la_data_in[23] la_data_out[18] la_data_in[96]
+ io_in_3v3[10] io_oeb[1] la_data_out[41] wbs_adr_i[3] la_data_out[35] la_oenb[28]
+ la_oenb[101] la_data_in[47] wbs_dat_i[31] la_oenb[75] gpio_analog[5] la_data_in[46]
+ io_analog[4] io_in_3v3[24] la_data_out[49] la_data_out[122] la_oenb[115] gpio_noesd[6]
+ gpio_analog[11] la_data_in[5] io_in[12] la_data_in[55] user_clock2 gpio_analog[2]
+ wbs_dat_o[7] wbs_sel_i[1] la_oenb[33] wbs_dat_i[13] la_data_out[80] la_data_out[4]
+ wbs_dat_o[6] io_in[21] la_data_in[109] vccd1 wbs_dat_o[1] gpio_analog[3] in_ring_0/vdda2
+ wbs_adr_i[19] la_data_in[10] io_analog[5] la_oenb[114] io_in_3v3[18] la_data_in[9]
+ la_data_in[108] la_data_out[126] la_oenb[73] wbs_adr_i[1] la_data_out[120] la_data_out[44]
+ la_data_in[26] la_oenb[113] la_oenb[14] la_data_out[84] la_data_in[114] io_out[0]
+ in_ring
.ends

