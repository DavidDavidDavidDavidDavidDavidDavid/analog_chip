* NGSPICE file created from padring_flat.ext - technology: sky130A

.subckt padring_flat
X0 a_41723_677112# in_ring_0/constant_gm_fingers_0.Vout a_43834_677960# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=4.3e+12p pd=3.172e+07u as=7.25e+12p ps=5.348e+07u w=5e+06u l=1e+06u
X1 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X2 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=3.235e+13p pd=2.2294e+08u as=1.3679e+14p ps=1.00302e+09u w=5e+06u l=500000u
R0 user_analog_project_wrapper_empty_0.vssd2 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_generic_m3 w=7.55e+07u l=1e+07u
X3 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X4 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=2.51e+13p pd=1.7004e+08u as=2.624e+14p ps=1.70496e+09u w=5e+06u l=150000u
X6 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=7.39e+13p pd=5.3956e+08u as=2.9e+13p ps=2.116e+08u w=5e+06u l=500000u
X7 a_24084_271906# a_24084_271906# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.25e+12p pd=5.348e+07u as=9.6e+12p ps=6.5e+07u w=2.5e+06u l=500000u
X8 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=2.075e+13p pd=1.383e+08u as=0p ps=0u w=5e+06u l=150000u
X9 a_287394_343809# in_ring_0/analog_mux_0.x16.B a_287588_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X10 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X11 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.17928e+14p pd=5.06904e+09u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=1e+06u
X12 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.304e+14p pd=8.5216e+08u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X13 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X14 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.82653e+14p ps=9.7052e+09u w=5e+06u l=150000u
X15 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.54e+13p ps=3.1816e+08u w=5e+06u l=500000u
X16 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X17 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X18 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X19 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X20 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X21 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X22 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# a_536916_284434# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X23 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X24 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X25 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X26 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X27 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X28 a_42819_684860# user_analog_project_wrapper_empty_0.io_analog[9] a_43026_690893# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=2.32e+13p pd=1.6928e+08u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X29 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.x5.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X30 user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=2.14535e+14p ps=1.68384e+09u w=5e+07u l=200000u
X31 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.595e+13p ps=1.1638e+08u w=5e+06u l=500000u
X32 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X33 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=1.595e+13p pd=1.1638e+08u as=0p ps=0u w=5e+06u l=500000u
X34 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540371_681998# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X35 a_287588_343809# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x8.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X36 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=2.555e+13p pd=1.8022e+08u as=0p ps=0u w=5e+06u l=1e+06u
X37 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X38 user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X39 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=1.595e+13p pd=1.1638e+08u as=0p ps=0u w=5e+06u l=500000u
X40 a_537154_685355# a_534722_685355# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X41 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X42 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X43 user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X44 a_287394_349409# in_ring_0/analog_mux_0.x2.B a_287588_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X45 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X46 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X47 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.83e+13p ps=1.2732e+08u w=5e+06u l=1e+06u
X48 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X49 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X50 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X51 a_287144_347009# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X52 a_534722_685355# a_537154_685355# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X53 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X54 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X55 user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=3.18606e+14p ps=2.87548e+09u w=5e+07u l=200000u
X56 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+13p ps=1.6928e+08u w=5e+06u l=1e+06u
X57 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X58 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+13p ps=5.2976e+08u w=5e+06u l=500000u
X59 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_287144_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X60 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X61 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X62 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X63 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X64 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X65 a_288390_347809# in_ring_0/analog_mux_0.x16.B a_288584_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X66 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X67 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X68 a_287588_349409# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x1.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X69 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X70 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X71 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X72 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.SIG9 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X73 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X74 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X75 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X76 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X77 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X78 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X79 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X80 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X81 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x2.A a_287588_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X82 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X83 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X84 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X85 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X86 a_287588_347809# in_ring_0/analog_mux_0.x2.B a_287394_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X87 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X88 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.74e+13p pd=1.2696e+08u as=0p ps=0u w=5e+06u l=1e+06u
X89 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X90 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X91 a_288584_347809# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X92 a_287394_345409# in_ring_0/analog_mux_0.x19.Y a_287144_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X93 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X94 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X95 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X96 user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X97 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X98 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X99 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X100 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X101 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=3.81686e+14p ps=3.65032e+09u w=5e+07u l=200000u
X102 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X103 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X104 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X105 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540371_681998# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X106 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X107 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# in_ring_0/analog_mux_0.SIG13 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X108 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X109 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X110 a_288390_343809# in_ring_0/analog_mux_0.x19.Y a_288140_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X111 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X112 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X113 a_42819_684860# user_analog_project_wrapper_empty_0.io_analog[8] a_40125_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X114 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.685e+13p ps=3.2874e+08u w=5e+06u l=500000u
X115 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X116 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X117 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X119 user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X120 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X121 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=1e+06u
R1 user_analog_project_wrapper_empty_0.vssa2 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_generic_m3 w=7.45e+07u l=2.6e+06u
X122 user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X123 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X124 user_analog_project_wrapper_empty_0.io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X125 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X126 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X127 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X128 a_287144_343809# in_ring_0/analog_mux_0.x19.A a_287394_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X129 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X130 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X131 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X133 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X134 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X136 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X137 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X138 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X139 in_ring_0/analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X140 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X141 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X142 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X143 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X144 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X145 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X146 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X147 a_288390_349409# in_ring_0/analog_mux_0.x19.A a_288140_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X148 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X149 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X150 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X151 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X152 in_ring_0/analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X153 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X154 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X155 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X156 a_17579_272227# user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.395e+13p ps=9.558e+07u w=5e+06u l=500000u
X157 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X158 user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X159 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X160 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X161 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X162 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X163 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_288140_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X164 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540916_680434# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X165 a_530722_289355# in_ring_0/analog_mux_0.SIG14 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X166 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X167 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X169 in_ring_0/analog_mux_0.x20.VPWR a_24084_271906# in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X170 a_287144_349409# in_ring_0/analog_mux_0.x19.Y a_287394_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X171 user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X172 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X173 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X174 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X175 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X176 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X177 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X178 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X179 user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X180 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X181 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X182 a_288140_347809# in_ring_0/analog_mux_0.x19.Y a_288390_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X183 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X184 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X185 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X187 a_288584_346209# in_ring_0/analog_mux_0.x2.B a_288390_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X188 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X189 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X190 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X191 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X192 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.SIG12 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X193 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X194 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X195 a_288140_344609# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X196 a_540916_680434# a_540371_681998# a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X197 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[1] a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.406e+07u as=0p ps=0u w=5e+06u l=500000u
X198 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X199 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X200 in_ring_0/analog_mux_0.SIG5 user_analog_project_wrapper_empty_0.gpio_analog[12] a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X201 user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X202 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X203 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X204 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X207 a_536916_284434# in_ring_0/analog_mux_0.SIG13 a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X208 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X209 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.x3.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X210 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X211 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# in_ring_0/analog_mux_0.SIG13 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X213 user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X214 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X215 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X216 in_ring_0/constant_gm_fingers_0.VDD a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X217 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+13p ps=4.232e+08u w=5e+06u l=500000u
X218 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X219 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X220 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X221 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X222 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x16.A a_288584_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X223 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X225 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.83e+13p pd=1.2732e+08u as=0p ps=0u w=5e+06u l=150000u
X226 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X227 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X228 user_analog_project_wrapper_empty_0.io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X229 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X230 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.SIG11 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X231 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X232 a_287144_348609# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X233 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X234 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X235 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X236 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.81686e+14p pd=3.65032e+09u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X237 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.105e+13p pd=7.674e+07u as=0p ps=0u w=1.25e+06u l=1e+06u
X238 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X239 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X240 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X241 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X242 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X243 a_17579_272227# user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X244 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X245 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X246 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X247 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X248 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X249 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X250 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X251 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X252 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X253 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X254 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X255 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x2.A a_287588_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X256 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X257 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X258 a_41723_677112# in_ring_0/constant_gm_fingers_0.Vout a_43834_677960# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X259 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X260 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X261 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X262 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X263 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X264 a_287394_345409# in_ring_0/analog_mux_0.x16.B a_287588_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X265 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X266 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X267 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X268 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X269 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X270 user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X271 a_17579_272227# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X272 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X273 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X274 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X275 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X276 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X277 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X278 user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X279 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_287144_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X280 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X281 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X282 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X283 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X284 a_288390_343809# in_ring_0/analog_mux_0.x2.B a_288584_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X285 user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X286 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X287 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X288 a_287588_345409# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x6.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X289 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X290 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X291 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X292 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X293 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.SIG14 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X294 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X295 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X296 in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.gpio_analog[1] a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X297 a_17579_272227# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X298 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X299 in_ring_0/analog_mux_0.x20.VPWR a_24084_271906# a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X300 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X301 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X302 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X303 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X304 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X305 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X306 a_287588_343809# in_ring_0/analog_mux_0.x16.B a_287394_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X307 a_17579_272227# user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X308 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X309 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X310 a_288584_343809# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X311 user_analog_project_wrapper_empty_0.io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X312 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X313 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_287144_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X314 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X315 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X317 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X318 user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.406e+07u as=0p ps=0u w=5e+06u l=1e+06u
X319 a_288390_349409# in_ring_0/analog_mux_0.x16.B a_288584_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X320 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X321 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X322 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X323 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X324 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X325 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X326 a_540459_681940# user_analog_project_wrapper_empty_0.io_analog[0] a_540271_687858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X327 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X328 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X329 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X330 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X331 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X332 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X333 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X334 in_ring_0/constant_gm_fingers_0.VSS a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X335 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_288140_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X336 a_43026_690893# user_analog_project_wrapper_empty_0.io_analog[9] a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X337 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X338 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X339 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X340 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X341 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X342 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X343 a_287588_349409# in_ring_0/analog_mux_0.x2.B a_287394_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X344 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X345 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X346 a_288584_349409# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X347 a_287394_347009# in_ring_0/analog_mux_0.x19.A a_287144_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X348 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X349 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X350 in_ring_0/constant_gm_fingers_0.VSS a_41723_677112# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X351 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X352 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X353 a_540916_680434# a_540916_680434# a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.348e+07u w=2.5e+06u l=500000u
X354 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X355 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X356 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X357 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X358 a_288584_347809# in_ring_0/analog_mux_0.x16.B a_288390_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X359 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X360 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X361 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 a_288390_345409# in_ring_0/analog_mux_0.x19.A a_288140_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X363 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X364 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X365 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X366 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X367 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X368 in_ring_0/constant_gm_fingers_0.Vout a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=4.35e+12p pd=3.174e+07u as=0p ps=0u w=5e+06u l=1e+06u
X369 a_29040_272091# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X370 in_ring_0/constant_gm_fingers_0.VDD a_43834_677960# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X371 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X372 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X373 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X374 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X375 in_ring_0/analog_mux_0.SIG6 a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X376 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X377 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X378 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X379 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X380 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X381 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X382 a_287144_345409# in_ring_0/analog_mux_0.x19.Y a_287394_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X383 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X384 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X385 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X386 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X387 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X388 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[1] a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X389 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X390 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X391 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X392 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X393 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X394 a_24084_271906# in_ring_0/analog_mux_0.SIG6 a_29040_272091# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X395 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X396 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X397 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X398 a_540459_681940# user_analog_project_wrapper_empty_0.io_analog[0] a_540271_687858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X399 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X400 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X401 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X402 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X403 a_288140_343809# in_ring_0/analog_mux_0.x19.Y a_288390_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X404 user_analog_project_wrapper_empty_0.io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X405 a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X406 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X407 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X408 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X409 a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[8] a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X410 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# in_ring_0/analog_mux_0.SIG13 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X411 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X412 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X413 user_analog_project_wrapper_empty_0.io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X414 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X415 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.SIG11 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X416 in_ring_0/analog_mux_0.SIG5 user_analog_project_wrapper_empty_0.gpio_analog[12] a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X417 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X418 a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[8] a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X419 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X420 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X421 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X422 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X424 a_17579_272227# user_analog_project_wrapper_empty_0.gpio_analog[13] a_14374_271026# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X425 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X426 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X427 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X428 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X429 a_536459_285940# user_analog_project_wrapper_empty_0.gpio_analog[0] a_536271_291858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X430 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X431 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X432 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X433 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X434 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.x8.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X435 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X436 a_288140_349409# in_ring_0/analog_mux_0.x19.A a_288390_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X437 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X438 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X439 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X440 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X441 in_ring_0/constant_gm_fingers_0.VSS a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X442 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X443 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X444 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X445 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X446 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X447 user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X448 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X449 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X450 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X451 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X452 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X453 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X454 in_ring_0/constant_gm_fingers_0.VSS a_41723_677112# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X455 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X456 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X457 a_288140_346209# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X458 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X459 a_287144_344609# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X460 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X461 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X462 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X463 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X464 a_42819_684860# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X465 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X466 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X467 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X468 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X469 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X470 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.x1.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X471 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540916_680434# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X472 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X473 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X474 user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X475 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X476 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X477 a_29040_272091# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X478 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X479 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X480 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X481 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X482 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X483 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X484 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X485 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x16.A a_288584_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X486 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X487 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X488 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x2.A a_287588_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X489 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X490 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X491 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X492 user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X493 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X494 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X495 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X496 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X497 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.SIG14 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X498 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X499 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X500 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X501 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X502 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X503 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X504 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X505 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X506 in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.gpio_analog[1] a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X507 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X508 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X509 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X510 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X511 a_536459_285940# user_analog_project_wrapper_empty_0.gpio_analog[0] a_536271_291858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X512 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X513 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X514 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X515 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X516 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X517 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X518 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X519 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X521 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X522 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X523 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X524 in_ring_0/constant_gm_fingers_0.VSS a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X525 a_24084_271906# a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X526 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X527 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X528 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X529 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X530 a_287394_348609# in_ring_0/analog_mux_0.x19.Y a_287144_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X531 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X532 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X533 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X534 a_287394_347009# in_ring_0/analog_mux_0.x2.B a_287588_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X535 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X536 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.SIG15 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X537 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X538 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X539 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X540 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X541 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X542 a_14374_271026# user_analog_project_wrapper_empty_0.gpio_analog[13] a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X543 in_ring_0/analog_mux_0.x20.VPWR a_24084_271906# in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X544 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X545 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X546 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X547 in_ring_0/constant_gm_fingers_0.Vout a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X548 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X549 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X550 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X551 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_287144_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X552 a_29040_272091# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X553 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X554 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X555 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X556 in_ring_0/constant_gm_fingers_0.Vout a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.4192e+12p pd=1.168e+07u as=0p ps=0u w=2.5e+06u l=500000u
X557 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X558 a_288390_345409# in_ring_0/analog_mux_0.x2.B a_288584_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X559 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X560 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X561 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.SIG15 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X562 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X563 a_42819_684860# user_analog_project_wrapper_empty_0.io_analog[8] a_40125_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X564 a_287588_347009# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x4.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X565 a_41723_677112# in_ring_0/constant_gm_fingers_0.Vout a_43834_677960# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X566 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X567 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X568 user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X569 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X570 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X571 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X572 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X573 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X574 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X575 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_288140_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X576 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X577 in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.gpio_analog[1] a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X578 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X579 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X580 a_287588_345409# in_ring_0/analog_mux_0.x16.B a_287394_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X581 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X582 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X583 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X584 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X585 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X586 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X587 a_288584_345409# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X588 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X589 a_42819_684860# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X590 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X591 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X592 user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X593 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X594 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X595 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X596 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X597 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X598 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X599 a_537154_685355# a_534722_685355# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X600 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X601 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X602 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X603 user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X604 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X605 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X606 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X607 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X608 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X609 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X610 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X611 a_288584_343809# in_ring_0/analog_mux_0.x2.B a_288390_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X612 user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X613 in_ring_0/analog_mux_0.SIG14 a_530722_289355# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X614 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X615 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X616 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X617 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X618 a_534722_685355# a_537154_685355# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X619 user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X620 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_288140_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X621 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540916_680434# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X622 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X623 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X624 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X625 user_analog_project_wrapper_empty_0.io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X626 user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X627 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X628 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X629 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X630 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X631 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X632 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X633 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X634 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X635 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X636 a_43834_677960# in_ring_0/constant_gm_fingers_0.Vout a_41723_677112# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X637 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X638 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X639 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X640 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X641 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X642 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X643 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X644 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X645 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X646 a_29040_272091# in_ring_0/analog_mux_0.SIG6 a_24084_271906# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X647 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X648 a_288584_349409# in_ring_0/analog_mux_0.x16.B a_288390_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X649 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X650 a_29040_272091# in_ring_0/analog_mux_0.SIG6 a_24084_271906# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X651 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X652 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X653 a_288390_347009# in_ring_0/analog_mux_0.x19.Y a_288140_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X654 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X655 a_540371_681998# a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X656 user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X657 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X658 a_288140_347809# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X659 a_540916_680434# a_540371_681998# a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X660 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X661 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X662 a_42819_684860# user_analog_project_wrapper_empty_0.io_analog[9] a_43026_690893# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X663 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X664 user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X665 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X666 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X667 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X668 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X669 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X670 a_287144_347009# in_ring_0/analog_mux_0.x19.A a_287394_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X671 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X672 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X673 a_42819_684860# user_analog_project_wrapper_empty_0.io_analog[9] a_43026_690893# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X674 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X675 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X676 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X677 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X678 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X679 a_17579_272227# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X680 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X681 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X682 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X683 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X684 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X685 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x16.A a_288584_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X686 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X687 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X688 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X689 a_288140_345409# in_ring_0/analog_mux_0.x19.A a_288390_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X690 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X691 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X692 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[1] a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X693 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X694 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X695 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X696 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X697 in_ring_0/analog_mux_0.SIG6 a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X698 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X699 user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X700 a_540459_681940# user_analog_project_wrapper_empty_0.io_analog[0] a_540271_687858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X701 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X702 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X703 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X704 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X705 in_ring_0/analog_mux_0.x20.VPWR a_24084_271906# a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X706 a_14374_271026# user_analog_project_wrapper_empty_0.gpio_analog[13] a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X707 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X708 in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.gpio_analog[1] a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X709 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X710 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X711 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X712 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X713 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X714 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X715 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X716 user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X717 user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X718 a_536459_285940# user_analog_project_wrapper_empty_0.gpio_analog[0] a_536271_291858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X719 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.x6.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X720 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X721 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.SIG12 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X722 user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X723 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X724 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X726 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540371_681998# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X727 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# a_536916_284434# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X728 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X729 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X730 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X731 a_287394_348609# in_ring_0/analog_mux_0.x2.B a_287588_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X732 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X733 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X734 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X735 a_287144_346209# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X736 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X737 a_17579_272227# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X738 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X739 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X740 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X741 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X742 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X743 a_42819_684860# user_analog_project_wrapper_empty_0.io_analog[8] a_40125_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X744 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X745 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X746 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X747 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X748 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X749 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X750 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X751 in_ring_0/analog_mux_0.SIG5 a_11871_265693# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X752 a_287588_348609# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x2.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X753 user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X754 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X755 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X756 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X757 a_17579_272227# user_analog_project_wrapper_empty_0.gpio_analog[13] a_14374_271026# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X758 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X759 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X760 a_11871_265693# in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X761 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X762 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X763 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x2.A a_287588_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
R2 in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.vssd1 sky130_fd_pr__res_generic_m3 w=7.7e+07u l=5e+06u
X764 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X765 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X766 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X768 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X769 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X770 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X771 a_287394_344609# in_ring_0/analog_mux_0.x19.A a_287144_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X772 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X773 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X774 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X775 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X776 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X777 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X778 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X779 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X780 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X781 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X782 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X783 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X784 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.SIG9 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X785 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X786 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X787 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 a_43834_677960# in_ring_0/constant_gm_fingers_0.Vout a_41723_677112# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X789 a_43026_690893# user_analog_project_wrapper_empty_0.io_analog[9] a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X790 a_14374_271026# user_analog_project_wrapper_empty_0.gpio_analog[13] a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X791 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X792 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X793 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X794 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X795 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X796 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# in_ring_0/analog_mux_0.SIG13 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X797 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X798 in_ring_0/analog_mux_0.SIG14 a_530722_289355# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X799 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X800 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X801 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X802 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X803 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X804 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X805 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X806 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X807 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X808 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X809 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X810 a_540459_681940# user_analog_project_wrapper_empty_0.io_analog[0] a_540271_687858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X811 a_37693_693523# a_40125_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X812 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X813 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X814 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X815 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_287144_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X817 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X818 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X819 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X820 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X821 a_288390_348609# in_ring_0/analog_mux_0.x19.A a_288140_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X822 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# in_ring_0/analog_mux_0.SIG13 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X823 a_288390_347009# in_ring_0/analog_mux_0.x16.B a_288584_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X824 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X825 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X826 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X827 user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X828 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X829 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X830 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X831 user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X832 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X833 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X834 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X835 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X836 a_24084_271906# a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X837 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_288140_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X838 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X839 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X840 a_287144_348609# in_ring_0/analog_mux_0.x19.Y a_287394_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X841 in_ring_0/constant_gm_fingers_0.VSS a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X842 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X843 a_287588_347009# in_ring_0/analog_mux_0.x2.B a_287394_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X844 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X845 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X846 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X847 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X848 a_288584_347009# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X849 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X850 a_42819_684860# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X851 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X852 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540916_680434# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X853 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X854 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X855 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X856 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X857 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X858 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X859 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X860 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X861 a_14374_271026# user_analog_project_wrapper_empty_0.gpio_analog[13] a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X862 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X863 a_288584_345409# in_ring_0/analog_mux_0.x2.B a_288390_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X864 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X865 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X866 user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X867 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X868 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X869 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X870 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X871 a_536916_284434# in_ring_0/analog_mux_0.SIG13 a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X872 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X873 a_288140_343809# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X874 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X875 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X876 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X877 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X878 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X879 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X880 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X881 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X882 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X883 a_540371_681998# a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X884 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X885 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X886 a_536916_284434# in_ring_0/analog_mux_0.SIG13 a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X887 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X888 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X889 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X890 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X891 user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X892 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X893 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X894 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X895 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X896 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X897 in_ring_0/constant_gm_fingers_0.VDD a_43834_677960# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X898 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.SIG12 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X899 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X900 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x16.A a_288584_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X901 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X902 a_43834_677960# in_ring_0/constant_gm_fingers_0.Vout a_41723_677112# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X903 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X904 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X905 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X906 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X907 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X908 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X909 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X910 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X911 a_288140_349409# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X912 a_287144_347809# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X913 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X914 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X915 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X916 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X917 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X918 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X919 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X920 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X921 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X922 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540916_680434# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X923 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# a_536916_284434# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X924 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X925 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X926 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X927 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X928 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X929 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X930 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X931 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X932 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X933 in_ring_0/analog_mux_0.SIG5 a_11871_265693# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X934 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X935 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X936 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X937 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x16.A a_288584_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X938 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X939 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x2.A a_287588_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X940 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X941 in_ring_0/constant_gm_fingers_0.VDD a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X942 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X943 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X944 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X945 a_288140_347009# in_ring_0/analog_mux_0.x19.Y a_288390_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X946 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X947 a_11871_265693# in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X948 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.SIG11 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X949 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X950 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X951 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X952 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X953 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X954 in_ring_0/analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X955 a_540916_680434# a_540371_681998# a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X956 user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X957 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X958 a_287394_344609# in_ring_0/analog_mux_0.x16.B a_287588_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X959 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X960 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X961 a_536916_284434# in_ring_0/analog_mux_0.SIG13 a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X962 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X963 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540371_681998# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X964 a_42819_684860# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X965 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X966 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X967 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X968 a_43026_690893# user_analog_project_wrapper_empty_0.io_analog[9] a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X969 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X970 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X971 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X972 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.x4.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X973 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X974 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X975 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X976 a_17579_272227# user_analog_project_wrapper_empty_0.gpio_analog[13] a_14374_271026# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X977 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X978 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X979 a_287588_344609# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x7.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X980 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X981 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X982 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.SIG9 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X983 a_42819_684860# user_analog_project_wrapper_empty_0.io_analog[8] a_40125_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X984 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X985 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X986 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X987 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X988 user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X989 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X990 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X991 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X992 user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X993 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X994 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X995 a_37693_693523# a_40125_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X996 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X997 in_ring_0/analog_mux_0.x20.VPWR a_24084_271906# in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X998 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X999 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1000 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_287144_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1001 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1002 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1003 user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1004 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1005 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1006 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1007 user_analog_project_wrapper_empty_0.io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1008 a_288390_348609# in_ring_0/analog_mux_0.x16.B a_288584_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X1009 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1010 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1011 a_42819_684860# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1012 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1013 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1014 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1015 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1016 user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1017 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1018 user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1019 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.SIG14 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1020 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1021 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1022 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1023 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1024 a_287588_348609# in_ring_0/analog_mux_0.x2.B a_287394_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1025 a_288584_348609# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1026 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1027 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# a_536916_284434# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1028 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1029 a_287394_346209# in_ring_0/analog_mux_0.x19.Y a_287144_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X1030 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1031 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1032 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1034 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1035 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1036 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1037 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1038 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1039 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1040 user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1041 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1042 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1043 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1045 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1046 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1047 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1048 a_288390_344609# in_ring_0/analog_mux_0.x19.Y a_288140_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X1049 in_ring_0/analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1050 user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1051 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1052 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1053 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1055 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1056 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1057 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1058 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1059 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1060 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R3 in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.vssa1 sky130_fd_pr__res_generic_m4 w=2.75e+07u l=2.8e+06u
X1061 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1062 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1063 a_17579_272227# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1064 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1065 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1066 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1067 a_287144_344609# in_ring_0/analog_mux_0.x19.A a_287394_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1068 a_540916_680434# a_540371_681998# a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1069 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1070 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[1] a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1071 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1072 user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1073 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1074 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1075 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1076 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1077 a_536916_284434# in_ring_0/analog_mux_0.SIG13 a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1078 a_540459_681940# user_analog_project_wrapper_empty_0.io_analog[0] a_540271_687858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1079 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1080 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1081 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1082 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1083 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1084 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1085 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1086 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1087 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1088 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1089 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1090 in_ring_0/constant_gm_fingers_0.Vout a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1091 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1092 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_288140_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1093 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1094 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1095 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1096 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1097 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1100 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1101 a_17579_272227# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1102 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1103 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1104 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1105 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1106 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1107 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1108 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1109 a_288140_348609# in_ring_0/analog_mux_0.x19.A a_288390_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1110 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1111 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1112 a_288584_347009# in_ring_0/analog_mux_0.x16.B a_288390_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1113 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1114 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1115 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1116 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1117 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1118 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1119 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1120 a_40125_693523# a_37693_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X1121 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1122 in_ring_0/analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1123 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1124 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1125 in_ring_0/analog_mux_0.SIG6 a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1126 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.SIG11 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1127 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1128 a_288140_345409# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1129 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1130 a_287144_343809# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1131 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1132 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1133 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1134 in_ring_0/analog_mux_0.x20.VPWR a_24084_271906# a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1135 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1136 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1137 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1138 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1139 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[1] a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1141 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1142 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.x2.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1143 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1144 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1145 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1146 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1147 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1148 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1149 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x16.A a_288584_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1150 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1151 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1152 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1153 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x2.A a_287588_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1154 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1155 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1156 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1157 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1158 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1159 a_287144_349409# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1160 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1161 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1162 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_5.Y in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1163 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1164 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1165 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1166 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1167 in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.gpio_analog[1] a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1168 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1169 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1170 in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1171 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1172 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1173 a_536459_285940# user_analog_project_wrapper_empty_0.gpio_analog[0] a_536271_291858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1174 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1175 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1176 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1177 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1178 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1179 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1180 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1181 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x2.A a_287588_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1182 user_analog_project_wrapper_empty_0.io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1183 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1184 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1185 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1186 a_43026_690893# user_analog_project_wrapper_empty_0.io_analog[9] a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1187 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1188 a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1189 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1190 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1191 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1192 a_287394_347809# in_ring_0/analog_mux_0.x19.A a_287144_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1193 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.Y in_ring_0/analog_mux_0.SIG14 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1194 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1195 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1196 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1197 a_287394_346209# in_ring_0/analog_mux_0.x16.B a_287588_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1198 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1199 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1200 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1201 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1202 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1203 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1204 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1205 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.vdda1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1206 user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1207 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1208 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1209 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[1] user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1210 in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X1211 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_287144_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1212 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1213 a_540916_680434# a_540916_680434# a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1214 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1215 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1216 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1217 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1218 a_288390_344609# in_ring_0/analog_mux_0.x2.B a_288584_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1219 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1220 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1221 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# a_536916_284434# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1222 in_ring_0/analog_mux_0.SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1223 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 a_536916_284434# a_536916_284434# in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1225 a_287588_346209# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x5.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1226 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1227 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1228 a_24084_271906# in_ring_0/analog_mux_0.SIG6 a_29040_272091# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1229 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1230 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1231 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1232 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1233 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1234 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1235 user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.io_analog[1] user_analog_project_wrapper_empty_0.vccd1 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1236 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1237 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1238 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1239 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1240 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1241 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1242 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1243 a_287588_344609# in_ring_0/analog_mux_0.x16.B a_287394_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1244 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1245 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1246 in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.gpio_analog[1] a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1247 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1248 a_288584_344609# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1249 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1250 user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1251 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1253 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1254 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1255 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.SIG15 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1256 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1257 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540371_681998# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1258 a_24084_271906# in_ring_0/analog_mux_0.SIG6 a_29040_272091# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1259 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1260 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1261 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1262 a_540459_681940# user_analog_project_wrapper_empty_0.io_analog[0] a_540271_687858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1263 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1264 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1265 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1266 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1267 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1268 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_288140_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1269 a_24084_271906# a_24084_271906# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1270 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1272 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1273 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1274 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1275 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1276 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1277 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1278 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1279 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1280 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1281 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1282 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1283 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1284 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1285 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 a_288584_348609# in_ring_0/analog_mux_0.x16.B a_288390_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1287 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1288 a_40125_693523# a_37693_693523# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X1289 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1290 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1291 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1292 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1293 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1294 a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1295 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1296 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1297 a_288390_346209# in_ring_0/analog_mux_0.x19.A a_288140_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1298 in_ring_0/constant_gm_fingers_0.VDD a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1299 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1300 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1301 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1302 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1303 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1304 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1305 user_analog_project_wrapper_empty_0.vdda1 user_analog_project_wrapper_empty_0.gpio_analog[0] user_analog_project_wrapper_empty_0.gpio_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1306 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1307 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1308 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1309 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_4.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1310 a_536916_284434# a_536916_284434# in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1311 user_analog_project_wrapper_empty_0.vccd1 user_analog_project_wrapper_empty_0.io_analog[0] user_analog_project_wrapper_empty_0.io_analog[0] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1312 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1313 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1314 a_287144_346209# in_ring_0/analog_mux_0.x19.Y a_287394_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1315 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1316 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1317 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1318 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1319 a_540371_681998# a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1320 user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1321 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1322 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1323 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1324 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1326 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1327 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1328 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1329 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1330 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1331 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1332 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1333 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1334 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1335 in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1336 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1337 in_ring_0/analog_mux_0.SIG6 a_24084_271906# a_24084_271906# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1338 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1339 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1340 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1341 a_288140_344609# in_ring_0/analog_mux_0.x19.Y a_288390_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1342 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1343 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1344 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1345 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1346 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1347 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1348 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1349 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1350 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1351 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1352 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1353 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1354 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1355 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1356 user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1357 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1358 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[13] user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1359 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1360 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1361 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1362 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1363 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1364 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1365 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1366 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1367 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1368 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1369 user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1370 user_analog_project_wrapper_empty_0.gpio_analog[13] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1371 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.x7.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1372 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1373 a_42819_684860# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1374 in_ring_0/constant_gm_fingers_0.VSS a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1375 a_536459_285940# user_analog_project_wrapper_empty_0.gpio_analog[0] a_536271_291858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1376 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1377 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1378 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1379 in_ring_0/analog_mux_0.SIG0 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1380 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1381 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1382 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1383 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1384 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1385 a_287394_347809# in_ring_0/analog_mux_0.x2.B a_287588_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1386 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1387 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1388 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1389 a_288140_347009# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1390 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1391 a_287144_345409# in_ring_0/analog_mux_0.x20.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1392 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1393 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540371_681998# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1394 user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1395 in_ring_0/analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1396 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1397 a_29040_272091# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X1398 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1399 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1400 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1401 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1402 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1403 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1404 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1405 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1406 a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[8] a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1407 in_ring_0/analog_mux_0.SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1408 a_29040_272091# in_ring_0/analog_mux_0.SIG6 a_24084_271906# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1409 a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1410 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1411 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1412 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1413 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1414 a_287588_347809# in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x3.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1415 a_40125_693523# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1416 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1417 user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1418 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1419 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1420 user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1421 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.A in_ring_0/analog_mux_0.x16.A a_288584_347009# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1422 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1423 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x2.A a_287588_345409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1424 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[1] a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1425 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1426 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.SIG1 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1427 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1428 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1429 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1430 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1431 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_3.Y in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1432 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1433 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1434 in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1435 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1436 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1437 a_287394_343809# in_ring_0/analog_mux_0.x19.A a_287144_343809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1438 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1439 in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.gpio_analog[1] a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1440 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1441 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1442 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.SIG15 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1443 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1444 in_ring_0/constant_gm_fingers_0.VSS a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1445 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1446 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1447 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1448 a_536459_285940# user_analog_project_wrapper_empty_0.gpio_analog[0] a_536271_291858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1449 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1450 in_ring_0/constant_gm_fingers_0.VSS a_41723_677112# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1451 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1452 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1453 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1454 a_540371_681998# a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1455 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1456 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1457 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1458 user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1459 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1460 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1461 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1463 in_ring_0/analog_mux_0.x1.Y in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1465 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.x2.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1466 user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1467 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1468 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1469 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1470 a_287394_349409# in_ring_0/analog_mux_0.x19.Y a_287144_349409# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1471 in_ring_0/analog_mux_0.SIG11 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1472 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1473 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1474 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1475 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1476 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1477 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1478 a_42819_684860# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1479 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1480 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1481 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1482 a_43834_677960# a_43834_677960# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1483 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1484 user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1485 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1486 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1487 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1488 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.Y in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1489 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1490 user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1491 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.SIG9 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1492 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.Y a_287144_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1493 in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X1494 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1495 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1496 a_288390_347809# in_ring_0/analog_mux_0.x19.Y a_288140_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1497 a_288390_346209# in_ring_0/analog_mux_0.x2.B a_288584_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1498 in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x16.B in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1499 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1500 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1501 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1502 in_ring_0/analog_mux_0.SIG5 user_analog_project_wrapper_empty_0.gpio_analog[12] a_17579_272227# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1503 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_1.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1504 user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1505 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.A a_288140_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1506 in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1507 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# in_ring_0/analog_mux_0.SIG13 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1508 a_540916_680434# a_540371_681998# a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1509 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1510 a_287144_347809# in_ring_0/analog_mux_0.x19.A a_287394_347809# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1511 in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1512 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1513 a_287588_346209# in_ring_0/analog_mux_0.x16.B a_287394_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1514 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1515 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1516 in_ring_0/analog_mux_0.SIG3 in_ring_0/analog_mux_0.x4.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1517 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 a_288584_346209# in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1519 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x16.B in_ring_0/analog_mux_0.x2.B in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1520 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1521 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1522 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1523 in_ring_0/analog_mux_0.SIG12 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1524 in_ring_0/analog_mux_0.x20.VPWR user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1525 user_analog_project_wrapper_empty_0.vccd1 a_540916_680434# a_540916_680434# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1526 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_2.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1528 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1529 a_540916_680434# a_540371_681998# a_541059_678436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1530 a_288584_344609# in_ring_0/analog_mux_0.x2.B a_288390_344609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1531 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1532 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1533 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1534 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1535 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1536 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1537 in_ring_0/constant_gm_fingers_0.VDD a_40125_693523# user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1538 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x16.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1539 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1540 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1541 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[1] a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1542 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_537154_685355# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1543 user_analog_project_wrapper_empty_0.gpio_analog[12] user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.x20.VPWR in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1544 in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_15.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1545 user_analog_project_wrapper_empty_0.io_analog[2] a_540371_681998# in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1546 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1547 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1548 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1549 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1550 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1551 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1552 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1553 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1554 in_ring_0/constant_gm_fingers_0.VSS a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X1555 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_6.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1556 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1557 in_ring_0/constant_gm_fingers_0.VSS a_41723_677112# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1558 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.A in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1559 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_43026_690893# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1560 a_540459_681940# user_analog_project_wrapper_empty_0.io_analog[0] a_540271_687858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1561 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# in_ring_0/analog_mux_0.SIG14 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1562 a_17579_272227# in_ring_0/analog_mux_0.SIG6 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1563 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1564 user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1565 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG13 a_536459_285940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1566 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout a_42819_684860# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1567 in_ring_0/constant_gm_fingers_0.VDD a_43026_690893# a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1568 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.gpio_analog[1] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1570 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1571 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_12.A in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1572 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x8.Y in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1573 a_536459_285940# user_analog_project_wrapper_empty_0.gpio_analog[0] a_536271_291858# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1574 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1575 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1576 a_530722_289355# in_ring_0/analog_mux_0.SIG14 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X1577 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.Y in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1578 in_ring_0/constant_gm_fingers_0.VSS a_540371_681998# a_540459_681940# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1579 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1580 in_ring_0/analog_mux_0.x20.VPWR a_14374_271026# in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1581 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1582 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1583 a_288140_348609# in_ring_0/analog_mux_0.x20.Y in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1584 user_analog_project_wrapper_empty_0.io_analog[10] a_40125_693523# in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1585 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x6.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1586 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_0.Y in_ring_0/analog_mux_0.SIG3 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1587 in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x19.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1588 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.Vout user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1589 in_ring_0/analog_mux_0.SIG5 a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1590 a_14374_271026# a_14374_271026# in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1591 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x3.Y in_ring_0/analog_mux_0.SIG2 in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1592 in_ring_0/analog_mux_0.SIG4 in_ring_0/analog_mux_0.x5.Y in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1593 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1594 in_ring_0/analog_mux_0.SIG7 in_ring_0/analog_mux_0.SIG5 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1595 user_analog_project_wrapper_empty_0.vdda1 in_ring_0/analog_mux_0.SIG14 in_ring_0/analog_mux_0.SIG15 user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1596 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1597 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_7.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1598 user_analog_project_wrapper_empty_0.io_analog[10] in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1599 in_ring_0/constant_gm_fingers_0.VSS a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X1600 in_ring_0/analog_mux_0.SIG15 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_14.A in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1601 in_ring_0/analog_mux_0.SIG9 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_8.Y in_ring_0/analog_mux_0.OUT in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1602 user_analog_project_wrapper_empty_0.vccd1 a_540271_687858# a_540271_687858# user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1603 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x19.A in_ring_0/analog_mux_0.x19.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1605 user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1606 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.A in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_10.A in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1607 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_9.A in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1608 in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.Y in_ring_0/analog_mux_0.x7.Y in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 in_ring_0/analog_mux_0.SIG13 in_ring_0/analog_mux_0.SIG13 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1610 in_ring_0/analog_mux_0.OUT in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_11.Y in_ring_0/analog_mux_0.SIG12 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1611 in_ring_0/analog_mux_0.sky130_fd_sc_hd__inv_2_13.A in_ring_0/analog_mux_0.x16.A a_288584_348609# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1612 in_ring_0/analog_mux_0.x2.Y in_ring_0/analog_mux_0.x2.B in_ring_0/analog_mux_0.x20.VPWR in_ring_0/analog_mux_0.x20.VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1613 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1614 user_analog_project_wrapper_empty_0.vdda1 a_536271_291858# a_536271_291858# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1615 user_analog_project_wrapper_empty_0.vdda1 a_536916_284434# a_536916_284434# user_analog_project_wrapper_empty_0.vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1616 in_ring_0/constant_gm_fingers_0.VDD user_analog_project_wrapper_empty_0.io_analog[8] user_analog_project_wrapper_empty_0.io_analog[8] in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1617 in_ring_0/constant_gm_fingers_0.VSS in_ring_0/analog_mux_0.SIG6 in_ring_0/analog_mux_0.SIG7 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1618 a_17579_272227# user_analog_project_wrapper_empty_0.gpio_analog[12] in_ring_0/analog_mux_0.SIG5 in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1619 a_288140_346209# in_ring_0/analog_mux_0.x19.A a_288390_346209# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1620 user_analog_project_wrapper_empty_0.io_analog[9] user_analog_project_wrapper_empty_0.io_analog[9] in_ring_0/constant_gm_fingers_0.VDD in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1621 user_analog_project_wrapper_empty_0.vccd1 a_537154_685355# user_analog_project_wrapper_empty_0.io_analog[2] user_analog_project_wrapper_empty_0.vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1622 a_536916_284434# in_ring_0/analog_mux_0.SIG13 a_537059_282436# in_ring_0/constant_gm_fingers_0.VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1623 in_ring_0/constant_gm_fingers_0.VDD a_43834_677960# in_ring_0/constant_gm_fingers_0.Vout in_ring_0/constant_gm_fingers_0.VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

