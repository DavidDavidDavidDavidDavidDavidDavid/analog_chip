** sch_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/user_analog_project_wrapper.sch
.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31]
+ wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23]
+ wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15]
+ wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7]
+ wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31]
+ wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28] wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23]
+ wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15]
+ wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[7]
+ wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24]
+ wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16]
+ wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8]
+ wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121]
+ la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114]
+ la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107]
+ la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100]
+ la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93]
+ la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79]
+ la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72]
+ la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58]
+ la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51]
+ la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44]
+ la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37]
+ la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30]
+ la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16]
+ la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9]
+ la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123]
+ la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117]
+ la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111]
+ la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98]
+ la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91]
+ la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77]
+ la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63]
+ la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56]
+ la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49]
+ la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42]
+ la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35]
+ la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28]
+ la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21]
+ la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14]
+ la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] io_in[26]
+ io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17] io_in[16] io_in[15]
+ io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4]
+ io_in[3] io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22]
+ io_in_3v3[21] io_in_3v3[20] io_in_3v3[19] io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14]
+ io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9] io_in_3v3[8] io_in_3v3[7] io_in_3v3[6]
+ io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] user_clock2 io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5]
+ io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22]
+ io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12]
+ io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13]
+ gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6]
+ gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] gpio_noesd[17]
+ gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10]
+ gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2]
+ gpio_noesd[1] gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5]
+ io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1]
+ io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_irq[2] user_irq[1] user_irq[0] la_oenb[127]
+ la_oenb[126] la_oenb[125] la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119]
+ la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111]
+ la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94]
+ la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85]
+ la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76]
+ la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69] la_oenb[68] la_oenb[67]
+ la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59] la_oenb[58]
+ la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49]
+ la_oenb[48] la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40]
+ la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31]
+ la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26] la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22]
+ la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13]
+ la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4]
+ la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0]
*.PININFO vdda1:B vdda2:B vssa1:B vssa2:B vccd1:B vccd2:B vssd1:B vssd2:B wb_clk_i:I wb_rst_i:I
*+ wbs_stb_i:I wbs_cyc_i:I wbs_we_i:I wbs_sel_i[3:0]:I wbs_dat_i[31:0]:I wbs_adr_i[31:0]:I wbs_ack_o:O
*+ wbs_dat_o[31:0]:O la_data_in[127:0]:I la_data_out[127:0]:O io_in[26:0]:I io_in_3v3[26:0]:I user_clock2:I
*+ io_out[26:0]:O io_oeb[26:0]:O gpio_analog[17:0]:B gpio_noesd[17:0]:B io_analog[10:0]:B io_clamp_high[2:0]:B
*+ io_clamp_low[2:0]:B user_irq[2:0]:O la_oenb[127:0]:I
XM2 net1 net5 net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=70 nf=14 m=1
XM1 net3 io_analog[9] net1 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM3 net4 io_analog[8] net1 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM4 net3 net3 vccd2 vccd2 sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM5 net4 net3 vccd2 vccd2 sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM6 io_analog[10] net4 vccd2 vccd2 sky130_fd_pr__pfet_01v8 L=0.5 W=200 nf=40 m=1
XM7 io_analog[10] net5 net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=60 nf=12 m=1
XC7 io_analog[10] net6 sky130_fd_pr__cap_mim_m3_1 W=16 L=16 MF=4 m=4
XR12 net6 net4 net2 sky130_fd_pr__res_xhigh_po_5p73 L=10 mult=4 m=4
XM8 net5 net7 vccd2 vccd2 sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM9 net7 net7 vccd2 vccd2 sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM10 net7 net5 net8 net2 sky130_fd_pr__nfet_01v8 L=1 W=30 nf=6 m=1
XM11 net5 net5 net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=4 m=1
XM12 net7 net7 net5 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=2 m=1
XR1 net2 net8 net2 sky130_fd_pr__res_xhigh_po_5p73 L=69 mult=4 m=4
XM13 net9 io_analog[0] net11 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=7
XM14 net11 net12 net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=14
XM15 net10 io_analog[1] net11 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=7
XM16 io_analog[2] net12 net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=12
XM17 net9 net9 vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=.5 W=5 nf=1 m=21
XM18 net10 net9 vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=.5 W=5 nf=1 m=21
XM19 io_analog[2] net10 vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=.5 W=5 nf=1 m=40
XR2 net15 net10 net2 sky130_fd_pr__res_xhigh_po_5p73 L=10 mult=4 m=4
XC1 io_analog[2] net15 sky130_fd_pr__cap_mim_m3_1 W=16 L=16 MF=4 m=4
XM33 net12 net13 vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 m=6
XM34 net13 net13 vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 m=6
XM35 net13 net12 net14 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=6
XM36 net12 net12 net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=1.25 nf=1 m=4
XM37 net13 net13 net12 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=2.5 nf=1 m=2
XR13 net2 net14 net2 sky130_fd_pr__res_xhigh_po_5p73 L=69 mult=4 m=4
R5 vssa1 net2 sky130_fd_pr__res_generic_m4 W=27.5 L=2.8 m=1
R4 vssa2 net2 sky130_fd_pr__res_generic_m3 W=74.5 L=2.6 m=1
XM20 net2 net2 io_analog[9] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM21 net2 net2 io_analog[8] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM22 io_analog[9] io_analog[9] vccd2 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM23 io_analog[8] io_analog[8] vccd2 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM24 net2 net2 io_analog[0] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM25 io_analog[0] io_analog[0] vccd1 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM26 net2 net2 io_analog[1] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM27 io_analog[1] io_analog[1] vccd1 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
x1 multiplier_vout multiplier_vmid multiplier_gm_voltage gpio_analog[16] gpio_analog[15] net2
+ gpio_analog[14] vdda2 fingers_vout fingers_gm_voltage fingers_vmid gpio_analog[11] gpio_analog[10] gpio_analog[9]
+ gpio_analog[8] gpio_analog[7] vdda2 net2 gpio_analog[6] gpio_analog[5] gpio_analog[4] gpio_analog[3]
+ gpio_analog[2] analog_mux
XM28 net16 fingers_gm_voltage net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=70 nf=14 m=1
XM29 net17 gpio_analog[13] net16 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM30 fingers_vmid gpio_analog[12] net16 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM31 net17 net17 vdda2 vdda2 sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM32 fingers_vmid net17 vdda2 vdda2 sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM38 fingers_vout fingers_vmid vdda2 vdda2 sky130_fd_pr__pfet_01v8 L=0.5 W=200 nf=40 m=1
XM39 fingers_vout fingers_gm_voltage net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=60 nf=12 m=1
XC2 fingers_vout net18 sky130_fd_pr__cap_mim_m3_1 W=16 L=16 MF=4 m=4
XR6 net18 fingers_vmid net2 sky130_fd_pr__res_xhigh_po_5p73 L=10 mult=4 m=4
XM40 fingers_gm_voltage net19 vdda2 vdda2 sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM41 net19 net19 vdda2 vdda2 sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM42 net19 fingers_gm_voltage net20 net2 sky130_fd_pr__nfet_01v8 L=1 W=30 nf=6 m=1
XM43 fingers_gm_voltage fingers_gm_voltage net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=4 m=1
XM44 net19 net19 fingers_gm_voltage net2 sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=2 m=1
XR8 net2 net20 net2 sky130_fd_pr__res_xhigh_po_5p73 L=69 mult=4 m=4
XM45 net21 gpio_analog[0] net22 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=7
XM46 net22 multiplier_gm_voltage net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=14
XM47 multiplier_vmid gpio_analog[1] net22 net2 sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=7
XM48 multiplier_vout multiplier_gm_voltage net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=12
XM49 net21 net21 vdda1 vdda1 sky130_fd_pr__pfet_01v8 L=.5 W=5 nf=1 m=21
XM50 multiplier_vmid net21 vdda1 vdda1 sky130_fd_pr__pfet_01v8 L=.5 W=5 nf=1 m=21
XM51 multiplier_vout multiplier_vmid vdda1 vdda1 sky130_fd_pr__pfet_01v8 L=.5 W=5 nf=1 m=40
XR10 net25 multiplier_vmid net2 sky130_fd_pr__res_xhigh_po_5p73 L=10 mult=4 m=4
XC3 multiplier_vout net25 sky130_fd_pr__cap_mim_m3_1 W=16 L=16 MF=4 m=4
XM52 multiplier_gm_voltage net23 vdda1 vdda1 sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 m=6
XM53 net23 net23 vdda1 vdda1 sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 m=6
XM54 net23 multiplier_gm_voltage net24 net2 sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=6
XM55 multiplier_gm_voltage multiplier_gm_voltage net2 net2 sky130_fd_pr__nfet_01v8 L=1 W=1.25 nf=1
+ m=4
XM56 net23 net23 multiplier_gm_voltage net2 sky130_fd_pr__nfet_01v8 L=0.5 W=2.5 nf=1 m=2
XR14 net2 net24 net2 sky130_fd_pr__res_xhigh_po_5p73 L=69 mult=4 m=4
R15 vssd1 net2 sky130_fd_pr__res_generic_m3 W=5 L=77 m=1
R16 vssd2 net2 sky130_fd_pr__res_generic_m3 W=10 L=75.5 m=1
XM57 net2 net2 gpio_analog[13] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM58 net2 net2 gpio_analog[12] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM59 gpio_analog[13] gpio_analog[13] vdda2 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM60 gpio_analog[12] gpio_analog[12] vdda2 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM61 net2 net2 gpio_analog[0] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM62 gpio_analog[0] gpio_analog[0] vdda1 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM63 net2 net2 gpio_analog[1] net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM64 gpio_analog[1] gpio_analog[1] vdda1 net2 sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
.ends

* expanding   symbol:  analog_mux.sym # of pins=23
** sym_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/analog_mux.sym
** sch_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/analog_mux.sch
.subckt analog_mux SIG15 SIG14 SIG13 SIG12 SIG11 SIG10 SIG9 SIG8 SIG7 SIG6 SIG5 SIG4 SIG3 SIG2 SIG1
+ SIG0 VDD GND SEL0 SEL1 SEL2 SEL3 OUT
*.PININFO OUT:O VDD:I GND:I SEL0:I SEL1:I SEL2:I SEL3:I SIG3:I SIG2:I SIG1:I SIG0:I SIG7:I SIG6:I
*+ SIG5:I SIG4:I SIG11:I SIG10:I SIG9:I SIG8:I SIG15:I SIG14:I SIG13:I SIG12:I
x1 VDD GND SEL0 SEL1 SEL2 SEL3 net1 net2 net4 net3 net5 net6 net8 net7 net9 net10 net12 net11 net13
+ net14 net16 net15 net17 net18 net20 net19 net21 net22 net24 net23 net25 net26 net28 net27 net29 net30
+ net32 net31 decoder_x4
x2 SIG15 net1 net2 SIG14 net4 net3 SIG13 net5 net6 SIG12 net8 net7 SIG11 net9 net10 SIG10 net12
+ net11 SIG9 net13 net14 SIG8 net16 net15 OUT SIG7 net17 net18 SIG6 net20 net19 SIG5 net21 net22 SIG4 net24
+ net23 SIG3 net25 net26 SIG2 net28 net27 SIG1 net29 net30 SIG0 net32 net31 VDD GND switch_x16
.ends


* expanding   symbol:  decoder_x4.sym # of pins=38
** sym_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/decoder_x4.sym
** sch_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/decoder_x4.sch
.subckt decoder_x4 VPWR VGND S0 S1 S2 S3 Q15N Q15 Q14N Q14 Q13N Q13 Q12N Q12 Q11N Q11 Q10N Q10 Q9N
+ Q9 Q8N Q8 Q7N Q7 Q6N Q6 Q5N Q5 Q4N Q4 Q3N Q3 Q2N Q2 Q1N Q1 Q0N Q0
*.PININFO S3:I S2:I S1:I S0:I VGND:I VPWR:I Q14N:O Q15N:O Q13N:O Q12N:O Q10N:O Q11N:O Q9N:O Q8N:O
*+ Q7N:O Q6N:O Q4N:O Q3N:O Q2N:O Q1N:O Q0N:O Q5N:O Q14:O Q15:O Q13:O Q12:O Q10:O Q11:O Q9:O Q8:O Q7:O Q6:O
*+ Q4:O Q3:O Q2:O Q1:O Q0:O Q5:O
x17 S3 VGND VGND VPWR VPWR S3N sky130_fd_sc_hd__inv_8
x18 S2 VGND VGND VPWR VPWR S2N sky130_fd_sc_hd__inv_8
x19 S1 VGND VGND VPWR VPWR S1N sky130_fd_sc_hd__inv_8
x20 S0 VGND VGND VPWR VPWR S0N sky130_fd_sc_hd__inv_8
x21 Q0N VGND VGND VPWR VPWR Q0 sky130_fd_sc_hd__inv_2
x22 Q1N VGND VGND VPWR VPWR Q1 sky130_fd_sc_hd__inv_2
x23 Q2N VGND VGND VPWR VPWR Q2 sky130_fd_sc_hd__inv_2
x24 Q3N VGND VGND VPWR VPWR Q3 sky130_fd_sc_hd__inv_2
x1 S3N S2N S1N S0N VGND VGND VPWR VPWR Q0N sky130_fd_sc_hd__nand4_2
x2 S3N S2N S1N S0 VGND VGND VPWR VPWR Q1N sky130_fd_sc_hd__nand4_2
x3 S3N S2N S1 S0N VGND VGND VPWR VPWR Q2N sky130_fd_sc_hd__nand4_2
x4 S3N S2N S1 S0 VGND VGND VPWR VPWR Q3N sky130_fd_sc_hd__nand4_2
x5 S3N S2 S1N S0N VGND VGND VPWR VPWR Q4N sky130_fd_sc_hd__nand4_2
x6 S3N S2 S1N S0 VGND VGND VPWR VPWR Q5N sky130_fd_sc_hd__nand4_2
x7 S3N S2 S1 S0N VGND VGND VPWR VPWR Q6N sky130_fd_sc_hd__nand4_2
x8 S3N S2 S1 S0 VGND VGND VPWR VPWR Q7N sky130_fd_sc_hd__nand4_2
x9 S3 S2N S1N S0N VGND VGND VPWR VPWR Q8N sky130_fd_sc_hd__nand4_2
x10 S3 S2N S1N S0 VGND VGND VPWR VPWR Q9N sky130_fd_sc_hd__nand4_2
x11 S3 S2N S1 S0N VGND VGND VPWR VPWR Q10N sky130_fd_sc_hd__nand4_2
x12 S3 S2N S1 S0 VGND VGND VPWR VPWR Q11N sky130_fd_sc_hd__nand4_2
x13 S3 S2 S1N S0N VGND VGND VPWR VPWR Q12N sky130_fd_sc_hd__nand4_2
x14 S3 S2 S1N S0 VGND VGND VPWR VPWR Q13N sky130_fd_sc_hd__nand4_2
x15 S3 S2 S1 S0N VGND VGND VPWR VPWR Q14N sky130_fd_sc_hd__nand4_2
x16 S3 S2 S1 S0 VGND VGND VPWR VPWR Q15N sky130_fd_sc_hd__nand4_2
x25 Q4N VGND VGND VPWR VPWR Q4 sky130_fd_sc_hd__inv_2
x26 Q5N VGND VGND VPWR VPWR Q5 sky130_fd_sc_hd__inv_2
x27 Q6N VGND VGND VPWR VPWR Q6 sky130_fd_sc_hd__inv_2
x28 Q7N VGND VGND VPWR VPWR Q7 sky130_fd_sc_hd__inv_2
x29 Q8N VGND VGND VPWR VPWR Q8 sky130_fd_sc_hd__inv_2
x30 Q9N VGND VGND VPWR VPWR Q9 sky130_fd_sc_hd__inv_2
x31 Q10N VGND VGND VPWR VPWR Q10 sky130_fd_sc_hd__inv_2
x32 Q11N VGND VGND VPWR VPWR Q11 sky130_fd_sc_hd__inv_2
x33 Q12N VGND VGND VPWR VPWR Q12 sky130_fd_sc_hd__inv_2
x34 Q13N VGND VGND VPWR VPWR Q13 sky130_fd_sc_hd__inv_2
x35 Q14N VGND VGND VPWR VPWR Q14 sky130_fd_sc_hd__inv_2
x36 Q15N VGND VGND VPWR VPWR Q15 sky130_fd_sc_hd__inv_2
.ends


* expanding   symbol:  switch_x16.sym # of pins=51
** sym_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/switch_x16.sym
** sch_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/switch_x16.sch
.subckt switch_x16 S15 PG15 NG15 S14 PG14 NG14 S13 PG13 NG13 S12 PG12 NG12 S11 PG11 NG11 S10 PG10
+ NG10 S9 PG9 NG9 S8 PG8 NG8 D S7 PG7 NG7 S6 PG6 NG6 S5 PG5 NG5 S4 PG4 NG4 S3 PG3 NG3 S2 PG2 NG2 S1 PG1
+ NG1 S0 PG0 NG0 VPB VNB
*.PININFO PG0:I NG0:I S0:I PG1:I NG1:I S1:I PG2:I NG2:I S2:I PG3:I NG3:I S3:I PG4:I NG4:I S4:I PG5:I
*+ NG5:I S5:I PG6:I NG6:I S6:I PG7:I NG7:I S7:I PG8:I NG8:I S8:I PG9:I NG9:I S9:I PG10:I NG10:I S10:I PG11:I
*+ NG11:I S11:I PG12:I NG12:I S12:I PG13:I NG13:I S13:I PG14:I NG14:I S14:I PG15:I NG15:I S15:I D:O VPB:I
*+ VNB:I
x1 S0 VNB NG0 VPB PG0 D a_mux_switch
x2 S1 VNB NG1 VPB PG1 D a_mux_switch
x3 S2 VNB NG2 VPB PG2 D a_mux_switch
x4 S3 VNB NG3 VPB PG3 D a_mux_switch
x5 S4 VNB NG4 VPB PG4 D a_mux_switch
x6 S5 VNB NG5 VPB PG5 D a_mux_switch
x7 S6 VNB NG6 VPB PG6 D a_mux_switch
x8 S7 VNB NG7 VPB PG7 D a_mux_switch
x9 S8 VNB NG8 VPB PG8 D a_mux_switch
x10 S9 VNB NG9 VPB PG9 D a_mux_switch
x11 S10 VNB NG10 VPB PG10 D a_mux_switch
x15 S11 VNB NG11 VPB PG11 D a_mux_switch
x16 S12 VNB NG12 VPB PG12 D a_mux_switch
x17 S13 VNB NG13 VPB PG13 D a_mux_switch
x18 S14 VNB NG14 VPB PG14 D a_mux_switch
x19 S15 VNB NG15 VPB PG15 D a_mux_switch
.ends


* expanding   symbol:  a_mux_switch.sym # of pins=6
** sym_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/a_mux_switch.sym
** sch_path: /foss/designs/C2S2_Analog_TestChip-main_3Outpus/xschem/a_mux_switch.sch
.subckt a_mux_switch VD VNB VNG VPB VPG VS
*.PININFO VPG:I VNG:I VD:I VS:O VPB:I VNB:I
XM1 VD VPG VS VPB sky130_fd_pr__pfet_01v8 L=0.15 W=95 nf=19 m=1
XM2 VD VNG VS VNB sky130_fd_pr__nfet_01v8 L=0.15 W=45 nf=9 m=1
.ends

.GLOBAL VPB
.GLOBAL VNB
.end
