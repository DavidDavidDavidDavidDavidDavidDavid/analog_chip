* NGSPICE file created from user_analog_project_wrapper_flat.ext - technology: sky130A

.subckt user_analog_project_wrapper_flat gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd2 vccd1 vdda2 vdda1
X0 a_41723_677112# a_42877_684772# a_43834_677960# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=4.3e+12p pd=3.172e+07u as=7.25e+12p ps=5.348e+07u w=5e+06u l=1e+06u
X1 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X2 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=3.235e+13p pd=2.2294e+08u as=1.3679e+14p ps=1.00302e+09u w=5e+06u l=500000u
R0 vssd2 a_5816_240836# sky130_fd_pr__res_generic_m3 w=7.55e+07u l=1e+07u
X3 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X4 a_286829_352328# a_284589_352318# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=2.51e+13p pd=1.7004e+08u as=2.624e+14p ps=1.70496e+09u w=5e+06u l=150000u
X6 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=7.39e+13p pd=5.3956e+08u as=2.9e+13p ps=2.116e+08u w=5e+06u l=500000u
X7 a_24084_271906# a_24084_271906# a_20532_271136# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=7.25e+12p pd=5.348e+07u as=9.6e+12p ps=6.5e+07u w=2.5e+06u l=500000u
X8 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=2.075e+13p pd=1.383e+08u as=0p ps=0u w=5e+06u l=150000u
X9 a_287394_343809# gpio_analog[4] a_287588_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X10 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X11 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=7.17928e+14p pd=5.06904e+09u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=1e+06u
X12 gpio_analog[2] a_284459_345646# gpio_analog[11] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.304e+14p pd=8.5216e+08u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X13 a_287812_343783# gpio_analog[3] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X14 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.82653e+14p ps=9.7052e+09u w=5e+06u l=150000u
X15 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.54e+13p ps=3.1816e+08u w=5e+06u l=500000u
X16 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X17 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X18 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X19 a_287139_344765# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X20 a_288222_346459# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X21 a_282219_342236# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X22 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X23 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X24 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X25 vdda2 a_287364_345383# a_288222_344059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X26 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X27 a_287139_344765# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X28 a_42819_684860# io_analog[9] a_43026_690893# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=2.32e+13p pd=1.6928e+08u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X29 a_284459_345646# a_282219_345636# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X30 io_analog[8] io_analog[8] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=2.14535e+14p ps=1.68384e+09u w=5e+07u l=200000u
X31 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.595e+13p ps=1.1638e+08u w=5e+06u l=500000u
X32 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X33 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=1.595e+13p pd=1.1638e+08u as=0p ps=0u w=5e+06u l=500000u
X34 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X35 a_287588_343809# a_287812_343783# a_284689_340388# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X36 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=2.555e+13p pd=1.8022e+08u as=0p ps=0u w=5e+06u l=1e+06u
X37 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X38 io_analog[8] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X39 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=1.595e+13p pd=1.1638e+08u as=0p ps=0u w=5e+06u l=500000u
X40 a_537154_685355# a_534722_685355# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X41 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X42 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X43 io_analog[9] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X44 a_287394_349409# a_287350_342628# a_287588_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X45 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X46 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X47 a_5816_240836# a_20532_271136# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.83e+13p ps=1.2732e+08u w=5e+06u l=1e+06u
X48 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X49 a_5816_240836# gpio_analog[6] a_287139_344765# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X50 a_5816_240836# gpio_analog[4] a_287350_342628# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X51 a_287144_347009# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X52 a_534722_685355# a_537154_685355# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X53 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X54 a_286876_343809# a_284689_340388# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X55 gpio_analog[13] gpio_analog[13] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=3.18606e+14p ps=2.87548e+09u w=5e+07u l=200000u
X56 a_5816_240836# a_20532_271136# a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+13p ps=1.6928e+08u w=5e+06u l=1e+06u
X57 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X58 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+13p ps=5.2976e+08u w=5e+06u l=500000u
X59 a_5816_240836# a_287139_344765# a_287144_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X60 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X61 a_5816_240836# a_42877_684772# a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X62 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X63 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X64 gpio_analog[7] a_286829_352328# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X65 a_288390_347809# gpio_analog[4] a_288584_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X66 a_282219_350736# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X67 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X68 a_287588_349409# a_287812_343783# a_284589_352318# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X69 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X70 a_289220_343809# a_288222_344059# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X71 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X72 gpio_analog[2] a_289220_344609# gpio_analog[14] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X73 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X74 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X75 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X76 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X77 a_20532_271136# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X78 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X79 vdda2 gpio_analog[13] gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X80 gpio_analog[16] a_289220_347009# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X81 a_282219_347336# a_287812_343783# a_287588_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X82 a_5816_240836# a_5816_240836# io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X83 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X84 a_282219_343936# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X85 vccd2 io_analog[9] io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X86 a_287588_347809# a_287350_342628# a_287394_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X87 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X88 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.74e+13p pd=1.2696e+08u as=0p ps=0u w=5e+06u l=1e+06u
X89 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X90 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X91 a_288584_347809# gpio_analog[3] a_288222_348059# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X92 a_287394_345409# a_287364_345383# a_287144_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X93 gpio_analog[2] a_284459_350746# gpio_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.15e+12p ps=5.326e+07u w=5e+06u l=150000u
X94 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X95 vdda2 a_287812_343783# a_282219_347336# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X96 gpio_analog[13] gpio_analog[13] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X97 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X98 gpio_analog[11] a_284459_345646# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X99 gpio_analog[16] a_289220_347009# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X100 a_288222_347259# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X101 io_analog[0] io_analog[0] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=3.81686e+14p ps=3.65032e+09u w=5e+07u l=200000u
X102 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X103 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X104 a_5816_240836# a_5816_240836# gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X105 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X106 a_289220_349409# a_288222_349659# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X107 vdda1 a_536916_284434# a_290737_348985# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X108 gpio_analog[11] a_284459_345646# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X109 gpio_analog[16] a_289220_347009# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X110 a_288390_343809# a_287364_345383# a_288140_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X111 a_287364_345383# gpio_analog[5] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X112 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X113 a_42819_684860# io_analog[8] a_40125_693523# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X114 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.685e+13p ps=3.2874e+08u w=5e+06u l=500000u
X115 vdda2 gpio_analog[3] a_288222_345659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X116 vccd2 io_analog[8] io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X117 vdda2 a_287350_342628# a_282219_347336# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 vccd1 io_analog[0] io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X119 io_analog[9] io_analog[9] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X120 a_5816_240836# a_42877_684772# a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X121 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=1e+06u
R1 vssa2 a_5816_240836# sky130_fd_pr__res_generic_m3 w=7.45e+07u l=2.6e+06u
X122 gpio_analog[12] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X123 a_5816_240836# a_5816_240836# io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X124 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X125 vdda2 gpio_analog[5] a_287364_345383# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X126 vdda2 gpio_analog[3] a_287812_343783# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X127 a_289220_347009# a_288222_347259# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X128 a_287144_343809# gpio_analog[5] a_287394_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X129 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X130 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X131 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 a_5816_240836# gpio_analog[5] a_287364_345383# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X133 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X134 vdda2 a_287350_342628# a_288222_345659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X136 io_analog[0] io_analog[0] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X137 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X138 a_288222_349659# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X139 a_12801_269626# a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X140 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X141 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X142 a_5816_240836# a_5816_240836# gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X143 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X144 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X145 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X146 a_5816_240836# a_288222_348059# a_289220_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X147 a_288390_349409# gpio_analog[5] a_288140_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X148 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X149 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X150 a_5816_240836# a_5816_240836# gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X151 gpio_analog[2] a_286829_352328# gpio_analog[7] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X152 a_12801_269626# a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X153 vdda2 a_282219_342236# a_284459_342246# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X154 gpio_analog[15] a_289220_346209# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X155 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X156 a_17579_272227# gpio_analog[12] a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.395e+13p ps=9.558e+07u w=5e+06u l=500000u
X157 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X158 io_analog[8] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X159 vccd1 io_analog[0] io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X160 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X161 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X162 a_287812_343783# gpio_analog[3] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X163 a_5816_240836# gpio_analog[6] a_288140_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X164 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X165 a_530722_289355# a_290737_350685# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X166 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X167 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 gpio_analog[12] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X169 vdda2 a_24084_271906# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X170 a_287144_349409# a_287364_345383# a_287394_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X171 gpio_analog[13] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X172 gpio_analog[2] a_286829_352328# gpio_analog[7] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X173 vdda2 a_288222_345659# a_289220_345409# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X174 a_288222_347259# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X175 a_5816_240836# a_5816_240836# io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X176 gpio_analog[8] a_284459_350746# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X177 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X178 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X179 gpio_analog[12] gpio_analog[12] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X180 io_analog[0] io_analog[0] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X181 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X182 a_288140_347809# a_287364_345383# a_288390_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X183 gpio_analog[8] a_284459_350746# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X184 a_5816_240836# a_5816_240836# gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X185 a_288222_344059# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X187 a_288584_346209# a_287350_342628# a_288390_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X188 a_5816_240836# gpio_analog[6] a_287139_344765# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X189 a_5816_240836# gpio_analog[4] a_287350_342628# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X190 vdda2 gpio_analog[5] a_282219_347336# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X191 gpio_analog[2] a_284459_345646# gpio_analog[11] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X192 gpio_analog[2] a_289220_347009# gpio_analog[16] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X193 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X194 vdda2 gpio_analog[13] gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X195 a_288140_344609# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X196 a_540916_680434# a_540371_681998# a_541059_678436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X197 a_537154_685355# io_analog[1] a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.406e+07u as=0p ps=0u w=5e+06u l=500000u
X198 a_5816_240836# a_282219_347336# a_284459_347346# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X199 a_287350_342628# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X200 a_11871_268125# gpio_analog[12] a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X201 gpio_analog[13] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X202 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X203 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X204 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 vdda2 gpio_analog[5] a_288222_345659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 gpio_analog[2] a_284459_345646# gpio_analog[11] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X207 a_536916_284434# a_290737_348985# a_537059_282436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X208 a_287350_342628# gpio_analog[4] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X209 a_284459_349046# a_282219_349036# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X210 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X211 vdda1 a_536916_284434# a_290737_348985# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X213 gpio_analog[13] gpio_analog[13] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X214 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X215 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X216 vccd2 a_43834_677960# a_43834_677960# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X217 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+13p ps=4.232e+08u w=5e+06u l=500000u
X218 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X219 a_12801_269626# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X220 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X221 a_5816_240836# a_5816_240836# gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X222 a_288222_344859# gpio_analog[3] a_288584_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X223 a_282219_342236# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X225 a_290737_350685# a_289220_348609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.83e+13p pd=1.2732e+08u as=0p ps=0u w=5e+06u l=150000u
X226 io_analog[1] io_analog[1] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X227 gpio_analog[7] a_286829_352328# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X228 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X229 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X230 gpio_analog[2] a_289220_346209# gpio_analog[15] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X231 a_5816_240836# a_42877_684772# a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X232 a_287144_348609# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X233 a_284459_343946# a_282219_343936# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X234 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X235 a_5816_240836# a_5816_240836# io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X236 vdda1 gpio_analog[1] gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.81686e+14p pd=3.65032e+09u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X237 a_290737_348985# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.105e+13p pd=7.674e+07u as=0p ps=0u w=1.25e+06u l=1e+06u
X238 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X239 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X240 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X241 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X242 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X243 a_17579_272227# gpio_analog[12] a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X244 gpio_analog[7] a_286829_352328# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X245 a_5816_240836# a_20532_271136# a_20532_271136# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X246 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X247 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X248 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X249 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X250 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X251 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X252 vdda2 gpio_analog[6] a_288222_348059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X253 vdda2 a_287139_344765# a_282219_345636# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X254 gpio_analog[7] a_286829_352328# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X255 a_282219_350736# a_287812_343783# a_287588_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X256 vccd1 io_analog[1] io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X257 gpio_analog[2] a_284459_350746# gpio_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X258 a_41723_677112# a_42877_684772# a_43834_677960# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X259 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X260 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X261 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X262 gpio_analog[1] gpio_analog[1] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X263 a_12801_269626# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X264 a_287394_345409# gpio_analog[4] a_287588_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X265 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X266 vdda2 gpio_analog[12] gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X267 vdda2 a_287812_343783# a_282219_350736# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X268 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X269 a_288222_348859# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X270 io_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X271 a_17579_272227# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X272 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X273 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X274 a_282219_345636# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X275 a_288222_348059# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X276 gpio_analog[2] a_284459_350746# gpio_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X277 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X278 gpio_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X279 a_5816_240836# gpio_analog[6] a_287144_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X280 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X281 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X282 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X283 a_287812_343783# gpio_analog[3] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X284 a_288390_343809# a_287350_342628# a_288584_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X285 gpio_analog[12] gpio_analog[12] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X286 a_282219_342236# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X287 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X288 a_287588_345409# a_287812_343783# a_282219_343936# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X289 vdda2 a_287350_342628# a_282219_350736# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X290 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.64e+13p ps=1.0656e+08u w=5e+06u l=150000u
X291 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X292 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X293 gpio_analog[2] a_289220_348609# a_290737_350685# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X294 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X295 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X296 a_290737_350685# gpio_analog[1] a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X297 a_17579_272227# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X298 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X299 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X300 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X301 gpio_analog[15] a_289220_346209# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X302 a_289220_348609# a_288222_348859# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X303 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X304 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X305 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X306 a_287588_343809# gpio_analog[4] a_287394_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X307 a_17579_272227# gpio_analog[12] a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X308 vdda2 gpio_analog[12] gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X309 a_5816_240836# gpio_analog[3] a_287812_343783# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X310 a_288584_343809# gpio_analog[3] a_288222_344059# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X311 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X312 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X313 a_5816_240836# a_287139_344765# a_287144_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X314 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X315 vdda2 gpio_analog[6] a_287139_344765# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X317 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X318 io_analog[10] a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.406e+07u as=0p ps=0u w=5e+06u l=1e+06u
X319 a_288390_349409# gpio_analog[4] a_288584_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X320 a_5816_240836# gpio_analog[6] a_287139_344765# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X321 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X322 gpio_analog[2] a_284459_343946# a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X323 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X324 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X325 gpio_analog[15] a_289220_346209# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X326 a_540459_681940# io_analog[0] a_540271_687858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X327 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X328 a_289220_345409# a_288222_345659# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X329 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X330 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X331 a_5816_240836# a_42877_684772# io_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X332 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X333 gpio_analog[2] a_286829_352328# gpio_analog[7] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X334 a_29040_272091# a_5816_240836# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.72e+06u l=6.9e+07u
X335 a_5816_240836# a_541059_678436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X336 a_5816_240836# gpio_analog[6] a_288140_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X337 a_43026_690893# io_analog[9] a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X338 gpio_analog[15] a_289220_346209# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X339 io_analog[1] io_analog[1] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X340 a_282219_347336# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X341 gpio_analog[9] a_284459_349046# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X342 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X343 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X344 a_287588_349409# a_287350_342628# a_287394_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X345 vdda2 a_289220_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X346 a_288222_348859# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X347 a_288584_349409# gpio_analog[3] a_288222_349659# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X348 a_287394_347009# gpio_analog[5] a_287144_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X349 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X350 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X351 a_5816_240836# a_41723_677112# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X352 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X353 vdda1 gpio_analog[1] gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X354 a_540916_680434# a_540916_680434# a_540371_681998# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.348e+07u w=2.5e+06u l=500000u
X355 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X356 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X357 a_288222_345659# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X358 gpio_analog[9] a_284459_349046# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X359 a_288584_347809# gpio_analog[4] a_288390_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X360 vdda2 a_287364_345383# a_282219_350736# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X361 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X362 a_5816_240836# a_288222_344059# a_289220_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X363 a_288390_345409# gpio_analog[5] a_288140_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X364 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X365 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X366 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=1.64e+13p pd=1.0656e+08u as=0p ps=0u w=5e+06u l=150000u
X367 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X368 vdda2 gpio_analog[3] a_288222_347259# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X369 a_42877_684772# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=4.35e+12p pd=3.174e+07u as=0p ps=0u w=5e+06u l=1e+06u
X370 vccd2 a_43834_677960# a_42877_684772# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X371 vccd1 io_analog[1] io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X372 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X373 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X374 a_5816_240836# a_289220_345409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X375 a_20532_271136# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X376 a_5816_240836# a_282219_350736# a_284459_350746# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X377 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X378 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X379 a_290737_350685# a_289220_348609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X380 gpio_analog[2] a_289220_347809# a_290737_348985# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X381 gpio_analog[1] gpio_analog[1] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X382 a_287144_345409# a_287364_345383# a_287394_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X383 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X384 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X385 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X386 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X387 vdda2 gpio_analog[4] a_288222_347259# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X388 a_537154_685355# io_analog[1] a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X389 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X390 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X391 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X392 a_5816_240836# a_288222_349659# a_289220_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X393 gpio_analog[2] a_286876_343809# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X394 a_24084_271906# a_20532_271136# a_29040_272091# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X395 a_290737_350685# a_289220_348609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X396 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X397 vdda2 a_282219_345636# a_284459_345646# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X398 a_540459_681940# io_analog[0] a_540271_687858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X399 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X400 a_11871_268125# a_284459_343946# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X401 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X402 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X403 a_288140_343809# a_287364_345383# a_288390_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X404 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X405 a_43834_677960# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X406 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X407 io_analog[0] io_analog[0] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X408 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X409 a_40125_693523# io_analog[8] a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X410 vdda1 a_536916_284434# a_290737_348985# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X411 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X412 a_290737_350685# a_289220_348609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X413 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X414 a_11871_268125# a_284459_343946# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X415 gpio_analog[2] a_289220_346209# gpio_analog[15] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X416 a_11871_268125# gpio_analog[12] a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X417 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X418 a_40125_693523# io_analog[8] a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X419 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X420 a_287364_345383# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X421 gpio_analog[2] a_289220_343809# vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X422 vdda2 a_288222_347259# a_289220_347009# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X424 a_17579_272227# gpio_analog[13] a_14374_271026# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X425 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X426 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X427 a_287364_345383# gpio_analog[5] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X428 vccd1 io_analog[0] io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X429 a_536459_285940# gpio_analog[0] a_536271_291858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X430 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X431 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X432 vdda2 gpio_analog[6] a_288222_349659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X433 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X434 a_286876_343809# a_284689_340388# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X435 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X436 a_288140_349409# gpio_analog[5] a_288390_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X437 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X438 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X439 gpio_analog[2] a_284459_349046# gpio_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X440 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X441 a_5816_240836# a_537059_282436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=6.9e+07u
X442 gpio_analog[2] a_289220_343809# vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X443 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X444 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X445 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X446 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X447 gpio_analog[13] gpio_analog[13] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X448 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X449 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X450 io_analog[0] io_analog[0] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X451 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X452 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X453 a_288447_352413# a_289220_349409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X454 a_5816_240836# a_41723_677112# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X455 a_5816_240836# gpio_analog[5] a_287364_345383# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X456 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X457 a_288140_346209# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X458 io_analog[1] io_analog[1] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X459 a_287144_344609# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X460 a_5816_240836# a_5816_240836# gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X461 gpio_analog[2] a_289220_345409# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X462 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X463 a_288222_349659# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X464 a_42819_684860# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X465 vdda2 a_287364_345383# a_288222_347259# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X466 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X467 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X468 a_5816_240836# a_20532_271136# a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X469 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X470 a_286829_352328# a_284589_352318# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X471 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X472 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X473 vdda2 gpio_analog[13] gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X474 io_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X475 vdda1 gpio_analog[0] gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X476 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X477 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X478 a_287139_344765# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X479 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X480 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X481 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X482 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X483 vdda2 a_287139_344765# a_288222_344059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X484 a_288222_346459# gpio_analog[3] a_288584_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X485 a_282219_345636# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X486 a_287139_344765# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X487 a_282219_342236# a_287812_343783# a_287588_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X488 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X489 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X490 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X491 gpio_analog[13] gpio_analog[13] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X492 a_5816_240836# a_20532_271136# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X493 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X494 a_284459_347346# a_282219_347336# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X495 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X496 gpio_analog[2] a_289220_348609# a_290737_350685# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X497 a_5816_240836# a_20532_271136# a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X498 a_290737_348985# a_289220_347809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X499 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X500 gpio_analog[2] a_284459_343946# a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X501 vdda2 a_287812_343783# a_282219_342236# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X502 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X503 a_288222_344859# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X504 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X505 a_290737_350685# gpio_analog[1] a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X506 a_5816_240836# a_5816_240836# io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X507 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X508 a_288222_344059# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X509 vdda2 gpio_analog[13] gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X510 a_536459_285940# gpio_analog[0] a_536271_291858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X511 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X512 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X513 a_12801_269626# a_286876_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X514 vdda2 a_287139_344765# a_282219_349036# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X515 gpio_analog[2] a_284459_343946# a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X516 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X517 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X518 vdda2 gpio_analog[4] a_282219_342236# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X519 a_282219_350736# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 gpio_analog[9] a_284459_349046# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X521 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X522 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X523 a_5816_240836# a_537059_282436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=6.9e+07u
X524 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X525 vdda2 a_289220_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X526 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X527 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X528 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X529 a_287394_348609# a_287364_345383# a_287144_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X530 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X531 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X532 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X533 a_287394_347009# a_287350_342628# a_287588_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X534 vdda2 gpio_analog[3] a_287812_343783# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X535 gpio_analog[2] a_289220_349409# a_288447_352413# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X536 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X537 a_289220_344609# a_288222_344859# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X538 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X539 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X540 vdda2 a_289220_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X541 a_14374_271026# gpio_analog[13] a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X542 vdda2 a_24084_271906# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X543 a_5816_240836# a_289220_345409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X544 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X545 a_282219_349036# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X546 a_42877_684772# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X547 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X548 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X549 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X550 a_5816_240836# gpio_analog[6] a_287144_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X551 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X552 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X553 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X554 a_42877_684772# a_43834_677960# a_43834_677960# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.4192e+12p pd=1.168e+07u as=0p ps=0u w=2.5e+06u l=500000u
X555 vccd1 io_analog[0] io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X556 a_288390_345409# a_287350_342628# a_288584_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X557 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X558 vdda2 gpio_analog[3] a_288222_348859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X559 gpio_analog[2] a_289220_349409# a_288447_352413# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X560 a_282219_345636# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X561 a_42819_684860# io_analog[8] a_40125_693523# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X562 a_287588_347009# a_287812_343783# a_282219_347336# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X563 a_41723_677112# a_42877_684772# a_43834_677960# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X564 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X565 gpio_analog[2] a_284459_342246# a_20532_271136# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X566 gpio_analog[13] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X567 a_5816_240836# a_289220_345409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X568 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X569 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X570 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X571 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X572 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X573 a_5816_240836# a_287139_344765# a_288140_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X575 a_290737_350685# gpio_analog[1] a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X576 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X577 a_5816_240836# a_289220_345409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X578 a_287588_345409# gpio_analog[4] a_287394_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X579 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X580 a_5816_240836# a_5816_240836# io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X581 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X582 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X583 a_288222_344859# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X584 vdda2 gpio_analog[4] a_288222_348859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X585 a_288584_345409# gpio_analog[3] a_288222_345659# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X586 gpio_analog[10] a_284459_347346# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=8.15e+12p pd=5.326e+07u as=0p ps=0u w=5e+06u l=150000u
X587 a_42819_684860# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X588 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X589 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X590 gpio_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X591 gpio_analog[2] a_289220_347809# a_290737_348985# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X592 a_5816_240836# a_5816_240836# gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X593 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X594 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X595 a_5816_240836# a_5816_240836# gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X596 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X597 a_537154_685355# a_534722_685355# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X598 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X599 vdda2 gpio_analog[4] a_287350_342628# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X600 a_5816_240836# a_42877_684772# a_42877_684772# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X601 io_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X602 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X603 a_5816_240836# gpio_analog[5] a_287364_345383# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X604 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X605 a_5816_240836# gpio_analog[3] a_287812_343783# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X606 a_289220_347009# a_288222_347259# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X607 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X608 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X609 a_288584_343809# a_287350_342628# a_288390_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X610 io_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X611 a_290737_350685# a_530722_289355# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X612 vdda2 gpio_analog[5] a_282219_342236# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X613 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X614 gpio_analog[2] a_286876_343809# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X615 gpio_analog[10] a_284459_347346# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X616 a_534722_685355# a_537154_685355# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X617 gpio_analog[13] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X618 a_5816_240836# gpio_analog[6] a_288140_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X619 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X620 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X621 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X622 a_12801_269626# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X623 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X624 gpio_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X625 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X626 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X627 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X628 vdda2 a_288222_348859# a_289220_348609# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X629 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X630 a_5816_240836# a_282219_342236# a_284459_342246# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X631 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X632 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X633 a_5816_240836# a_5816_240836# gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X634 a_43834_677960# a_42877_684772# a_41723_677112# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X635 a_5816_240836# a_5816_240836# io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X636 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X637 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X638 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X639 gpio_analog[2] a_289220_343809# vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X640 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X641 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X642 a_5816_240836# a_5816_240836# gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X643 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X644 a_29040_272091# a_20532_271136# a_24084_271906# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X645 a_288222_347259# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X646 a_288584_349409# gpio_analog[4] a_288390_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X647 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X648 a_29040_272091# a_20532_271136# a_24084_271906# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X649 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X650 a_5816_240836# a_288222_345659# a_289220_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X651 a_288390_347009# a_287364_345383# a_288140_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X652 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X653 a_540371_681998# a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X654 io_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X655 a_288447_352413# a_289220_349409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X656 a_288140_347809# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X657 a_540916_680434# a_540371_681998# a_541059_678436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X658 a_20532_271136# a_284459_342246# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X659 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X660 a_42819_684860# io_analog[9] a_43026_690893# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X661 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X662 gpio_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X663 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X664 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X665 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X666 vdda2 gpio_analog[5] a_288222_348859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X667 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X668 a_287144_347009# gpio_analog[5] a_287394_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X669 vccd2 io_analog[9] io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X670 a_20532_271136# a_284459_342246# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X671 a_42819_684860# io_analog[9] a_43026_690893# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X672 gpio_analog[2] a_289220_345409# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X673 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X674 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X675 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X676 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X677 a_17579_272227# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X678 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X679 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X680 vdda2 a_287139_344765# a_288222_345659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X681 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X682 a_12801_269626# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X683 a_288222_348059# gpio_analog[3] a_288584_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X684 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X685 a_287350_342628# gpio_analog[4] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X686 vdda2 a_282219_349036# a_284459_349046# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X687 a_288140_345409# gpio_analog[5] a_288390_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X688 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X689 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X690 a_537154_685355# io_analog[1] a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X691 a_284459_350746# a_282219_350736# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X692 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X693 gpio_analog[2] a_284459_347346# gpio_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X694 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X695 a_20532_271136# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X696 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X697 io_analog[10] a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X698 a_540459_681940# io_analog[0] a_540271_687858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X699 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X700 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X701 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X702 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X703 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X704 a_14374_271026# gpio_analog[13] a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X705 a_5816_240836# a_5816_240836# io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X706 a_290737_350685# gpio_analog[1] a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X707 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X708 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X709 a_288222_345659# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X710 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X711 a_5816_240836# a_5816_240836# gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X712 a_287812_343783# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X713 gpio_analog[14] a_289220_344609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X714 gpio_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X715 io_analog[10] a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X716 a_536459_285940# gpio_analog[0] a_536271_291858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X717 a_284459_343946# a_282219_343936# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X718 vdda2 a_287139_344765# a_284589_352318# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X719 gpio_analog[2] a_289220_347009# gpio_analog[16] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X720 io_analog[9] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X721 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X722 a_287139_344765# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X723 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X724 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X725 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X726 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X727 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X728 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X729 a_287394_348609# a_287350_342628# a_287588_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X730 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X731 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X732 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X733 a_287144_346209# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X734 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X735 a_17579_272227# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X736 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X737 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X738 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X739 a_284589_352318# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X740 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X741 a_42819_684860# io_analog[8] a_40125_693523# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X742 gpio_analog[2] a_284459_342246# a_20532_271136# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X743 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X744 a_5816_240836# a_5816_240836# io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X745 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X746 a_5816_240836# a_5816_240836# io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X747 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X748 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X749 a_11871_268125# a_11871_265693# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X750 a_287588_348609# a_287812_343783# a_282219_350736# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X751 io_analog[8] io_analog[8] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X752 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X753 vccd2 io_analog[9] io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X754 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X755 a_17579_272227# gpio_analog[13] a_14374_271026# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X756 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X757 a_5816_240836# a_5816_240836# gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X758 a_11871_265693# a_11871_268125# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X759 vdda2 gpio_analog[6] a_284689_340388# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X760 a_282219_349036# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X761 a_282219_345636# a_287812_343783# a_287588_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
R2 a_5816_240836# vssd1 sky130_fd_pr__res_generic_m3 w=7.7e+07u l=5e+06u
X762 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X763 gpio_analog[2] a_284459_342246# a_20532_271136# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X764 a_282219_342236# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X765 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X766 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X767 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X768 gpio_analog[10] a_284459_347346# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X769 a_287394_344609# gpio_analog[5] a_287144_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X770 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X771 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X772 vdda2 a_287812_343783# a_282219_345636# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X773 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X774 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X775 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X776 a_288222_346459# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X777 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X778 a_284689_340388# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X779 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X780 vccd2 io_analog[8] io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X781 a_289220_348609# a_288222_348859# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X782 gpio_analog[2] a_289220_344609# gpio_analog[14] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X783 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X784 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X785 vdda2 gpio_analog[3] a_288222_344859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X786 a_43834_677960# a_42877_684772# a_41723_677112# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X787 a_43026_690893# io_analog[9] a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X788 a_14374_271026# gpio_analog[13] a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X789 vdda2 gpio_analog[4] a_282219_345636# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X790 a_5816_240836# gpio_analog[6] a_287139_344765# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X791 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X792 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X793 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X794 vdda1 a_536916_284434# a_290737_348985# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X795 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X796 a_290737_350685# a_530722_289355# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X797 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X798 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X799 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X800 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X801 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X802 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X803 a_289220_346209# a_288222_346459# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X804 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X805 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X806 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X807 a_290737_348985# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X808 a_540459_681940# io_analog[0] a_540271_687858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X809 a_37693_693523# a_40125_693523# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X810 vdda2 a_287350_342628# a_288222_344859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X811 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X812 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X813 a_288222_348859# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X814 a_5816_240836# gpio_analog[6] a_287144_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X815 gpio_analog[11] a_284459_345646# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X816 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X817 gpio_analog[16] a_289220_347009# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X818 vdda2 gpio_analog[5] a_287364_345383# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X819 a_288390_348609# gpio_analog[5] a_288140_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X820 vdda1 a_536916_284434# a_290737_348985# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X821 a_288390_347009# gpio_analog[4] a_288584_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X822 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X823 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X824 a_282219_349036# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X825 io_analog[9] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X826 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X827 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X828 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X829 io_analog[9] io_analog[9] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X830 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X831 a_5816_240836# a_20532_271136# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X832 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X833 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X834 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X835 a_5816_240836# a_287139_344765# a_288140_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X836 gpio_analog[11] a_284459_345646# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X837 a_5816_240836# a_20532_271136# a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X838 a_287144_348609# a_287364_345383# a_287394_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X839 a_5816_240836# a_541059_678436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X840 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X841 a_287588_347009# a_287350_342628# a_287394_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X842 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X843 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X844 vdda2 a_288222_344859# a_289220_344609# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X845 a_288222_346459# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X846 a_288584_347009# gpio_analog[3] a_288222_347259# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X847 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X848 a_42819_684860# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X849 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X850 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X851 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X852 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X853 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X854 vdda2 a_284589_352318# a_286829_352328# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X855 a_5816_240836# a_42877_684772# io_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X856 gpio_analog[0] gpio_analog[0] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X857 a_20532_271136# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X858 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X859 a_14374_271026# gpio_analog[13] a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X860 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X861 a_288584_345409# a_287350_342628# a_288390_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X862 gpio_analog[14] a_289220_344609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X863 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X864 io_analog[8] io_analog[8] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X865 vdda2 a_287364_345383# a_282219_345636# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X866 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X867 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X868 vccd2 io_analog[9] io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X869 a_536916_284434# a_290737_348985# a_537059_282436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X870 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X871 a_288140_343809# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X872 a_5816_240836# a_42877_684772# a_42877_684772# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X873 vdda1 gpio_analog[0] gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X874 a_5816_240836# a_282219_345636# a_284459_345646# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X875 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X876 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X877 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X878 gpio_analog[14] a_289220_344609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X879 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X880 vdda2 a_287364_345383# a_288222_344859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X881 a_540371_681998# a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X882 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X883 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X884 a_536916_284434# a_290737_348985# a_537059_282436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X885 gpio_analog[14] a_289220_344609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X886 gpio_analog[8] a_284459_350746# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X887 a_287350_342628# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X888 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X889 io_analog[8] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X890 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X891 vccd2 io_analog[8] io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X892 gpio_analog[0] gpio_analog[0] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X893 a_287364_345383# gpio_analog[5] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X894 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X895 vccd2 a_43834_677960# a_42877_684772# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X896 gpio_analog[2] a_289220_347009# gpio_analog[16] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X897 a_5816_240836# a_288222_347259# a_289220_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X898 a_288222_344059# gpio_analog[3] a_288584_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X899 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X900 a_43834_677960# a_42877_684772# a_41723_677112# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X901 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X902 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X903 vdda2 a_284689_340388# a_286876_343809# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X904 a_5816_240836# a_5816_240836# io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X905 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X906 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X907 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X908 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X909 a_288140_349409# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X910 a_287144_347809# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X911 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X912 a_284459_342246# a_282219_342236# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X913 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X914 gpio_analog[8] a_284459_350746# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X915 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X916 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X917 vdda1 gpio_analog[0] gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X918 gpio_analog[2] a_284459_345646# gpio_analog[11] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X919 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X920 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X921 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X922 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X923 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X924 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X925 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X926 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X927 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X928 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X929 a_29040_272091# a_5816_240836# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.72e+06u l=6.9e+07u
X930 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X931 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X932 a_11871_268125# a_11871_265693# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X933 vdda2 a_287139_344765# a_288222_347259# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X934 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X935 vdda2 gpio_analog[6] a_282219_343936# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X936 a_288222_349659# gpio_analog[3] a_288584_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X937 a_284589_352318# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X938 a_282219_349036# a_287812_343783# a_287588_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X939 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X940 vccd2 a_43834_677960# a_43834_677960# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X941 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X942 gpio_analog[0] gpio_analog[0] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X943 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X944 a_288140_347009# a_287364_345383# a_288390_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X945 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X946 a_11871_265693# a_11871_268125# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X947 gpio_analog[2] a_289220_346209# gpio_analog[15] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X948 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X949 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X950 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X951 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X952 vccd2 io_analog[8] io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X953 a_288447_352413# a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X954 a_540916_680434# a_540371_681998# a_541059_678436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X955 io_analog[9] io_analog[9] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X956 a_287139_344765# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X957 a_287394_344609# gpio_analog[4] a_287588_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X958 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X959 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X960 a_536916_284434# a_290737_348985# a_537059_282436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X961 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X962 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X963 a_42819_684860# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X964 a_282219_343936# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X965 a_288222_347259# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X966 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X967 a_43026_690893# io_analog[9] a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X968 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X969 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X970 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X971 a_284459_347346# a_282219_347336# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X972 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X973 gpio_analog[7] a_286829_352328# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X974 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X975 a_17579_272227# gpio_analog[13] a_14374_271026# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X976 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X977 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X978 a_287588_344609# a_287812_343783# a_282219_342236# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X979 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X980 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X981 gpio_analog[2] a_289220_344609# gpio_analog[14] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X982 a_42819_684860# io_analog[8] a_40125_693523# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X983 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X984 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X985 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X986 a_5816_240836# a_5816_240836# io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X987 io_analog[8] io_analog[8] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X988 a_284689_340388# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X989 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X990 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X991 io_analog[8] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X992 gpio_analog[1] gpio_analog[1] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X993 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X994 a_37693_693523# a_40125_693523# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X995 a_5816_240836# a_5816_240836# gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X996 vdda2 a_24084_271906# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X997 gpio_analog[2] a_284459_350746# gpio_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X998 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X999 a_5816_240836# gpio_analog[6] a_287144_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1000 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1001 gpio_analog[11] a_284459_345646# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1002 io_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1003 vdda2 gpio_analog[3] a_287812_343783# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1004 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1005 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1006 io_analog[10] a_37693_693523# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1007 a_288390_348609# gpio_analog[4] a_288584_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.915e+11p ps=5.72e+06u w=650000u l=150000u
X1008 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1009 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1010 a_42819_684860# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1011 a_284589_352318# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1012 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1013 a_5816_240836# gpio_analog[3] a_287812_343783# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1014 a_289220_344609# a_288222_344859# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1015 gpio_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1016 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1017 gpio_analog[12] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1018 gpio_analog[2] a_289220_348609# a_290737_350685# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1019 a_5816_240836# a_5816_240836# io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1020 vdda1 gpio_analog[1] gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1021 a_5816_240836# a_5816_240836# io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1022 a_282219_345636# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1023 a_287588_348609# a_287350_342628# a_287394_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1024 a_288584_348609# gpio_analog[3] a_288222_348859# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1025 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1026 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1027 a_29040_272091# a_5816_240836# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.72e+06u l=6.9e+07u
X1028 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1029 a_287394_346209# a_287364_345383# a_287144_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X1030 a_5816_240836# a_5816_240836# gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1031 a_287350_342628# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1032 vdda2 a_287812_343783# a_282219_349036# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1034 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1035 a_288222_348059# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1036 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1037 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1038 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1039 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1040 io_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1041 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1042 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1043 a_288222_344859# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1045 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1046 a_5816_240836# a_42877_684772# io_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1047 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1048 a_288390_344609# a_287364_345383# a_288140_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X1049 a_288447_352413# a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1050 gpio_analog[0] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1051 gpio_analog[2] a_286829_352328# gpio_analog[7] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1052 vdda2 gpio_analog[3] a_288222_346459# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1053 vdda2 gpio_analog[4] a_287350_342628# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 gpio_analog[15] a_289220_346209# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1055 a_12801_269626# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1056 a_284689_340388# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1057 vdda2 a_287350_342628# a_282219_349036# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1058 a_5816_240836# a_42877_684772# io_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1059 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1060 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R3 a_5816_240836# vssa1 sky130_fd_pr__res_generic_m4 w=2.75e+07u l=2.8e+06u
X1061 a_5816_240836# gpio_analog[4] a_287350_342628# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1062 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1063 a_17579_272227# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1064 a_5816_240836# a_282219_349036# a_284459_349046# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1065 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1066 a_289220_347809# a_288222_348059# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1067 a_287144_344609# gpio_analog[5] a_287394_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1068 a_540916_680434# a_540371_681998# a_541059_678436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1069 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1070 a_537154_685355# io_analog[1] a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1071 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1072 io_analog[8] io_analog[8] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1073 vdda2 a_287350_342628# a_288222_346459# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1074 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1075 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1076 gpio_analog[8] a_284459_350746# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1077 a_536916_284434# a_290737_348985# a_537059_282436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1078 a_540459_681940# io_analog[0] a_540271_687858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1079 a_5816_240836# a_20532_271136# a_20532_271136# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1080 a_5816_240836# a_288222_348859# a_289220_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1081 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1082 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1083 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1084 vdda2 a_282219_343936# a_284459_343946# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1085 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1086 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1087 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1088 vdda2 gpio_analog[12] gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1089 vccd1 io_analog[1] io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1090 a_42877_684772# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1091 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1092 a_5816_240836# a_287139_344765# a_288140_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1093 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1094 a_29040_272091# a_5816_240836# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.72e+06u l=6.9e+07u
X1095 gpio_analog[1] gpio_analog[1] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1096 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1097 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1098 vdda2 a_288222_346459# a_289220_346209# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 a_288222_348059# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1100 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1101 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1102 a_17579_272227# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1103 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1104 vdda2 a_287139_344765# a_288222_348859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1105 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1106 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1107 vccd1 io_analog[1] io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1108 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1109 a_287364_345383# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1110 a_288140_348609# gpio_analog[5] a_288390_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1111 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1112 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1113 a_288584_347009# gpio_analog[4] a_288390_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1114 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1115 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1116 vdda2 gpio_analog[5] a_282219_349036# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1117 io_analog[1] io_analog[1] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1118 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1119 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1120 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1121 a_40125_693523# a_37693_693523# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X1122 a_290737_350685# a_289220_348609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1123 a_288447_352413# a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1124 gpio_analog[14] a_288222_344859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1125 a_11871_268125# a_284459_343946# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1126 a_20532_271136# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1127 gpio_analog[2] a_289220_346209# gpio_analog[15] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1128 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1129 a_288140_345409# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1130 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1131 a_287144_343809# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1132 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1133 a_5816_240836# a_42877_684772# a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1134 vdda1 gpio_analog[1] gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1135 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1136 a_288222_348859# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1137 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1138 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1139 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1140 vdda2 gpio_analog[5] a_288222_346459# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1141 a_537154_685355# io_analog[1] a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1142 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1143 a_284459_350746# a_282219_350736# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1144 a_11871_268125# a_284459_343946# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1145 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1146 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1147 gpio_analog[2] a_284459_349046# gpio_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1148 gpio_analog[2] a_288222_347259# gpio_analog[16] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1149 a_287812_343783# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1150 a_288222_345659# gpio_analog[3] a_288584_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1151 a_282219_343936# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1152 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1153 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1154 a_284689_340388# a_287812_343783# a_287588_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1155 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1156 a_287812_343783# gpio_analog[3] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1157 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1158 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1159 a_288447_352413# a_289220_349409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1160 a_287144_349409# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1161 a_287139_344765# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1162 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1163 a_284459_345646# a_282219_345636# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1164 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1165 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1166 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1167 gpio_analog[2] a_289220_345409# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1168 a_290737_350685# gpio_analog[1] a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1169 gpio_analog[0] gpio_analog[0] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1170 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1171 a_287139_344765# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1172 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1173 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1174 a_536459_285940# gpio_analog[0] a_536271_291858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1175 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1176 vdda2 gpio_analog[6] a_287139_344765# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1177 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1178 vdda2 gpio_analog[6] a_282219_347336# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1179 vdda2 gpio_analog[4] a_287350_342628# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1180 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1181 vdda1 gpio_analog[0] gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1182 a_284589_352318# a_287812_343783# a_287588_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1183 io_analog[2] a_534722_685355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1184 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1185 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1186 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1187 a_43026_690893# io_analog[9] a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1188 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1189 a_43834_677960# a_43834_677960# a_42877_684772# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1190 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1191 vccd1 io_analog[1] io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1192 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1193 a_287394_347809# gpio_analog[5] a_287144_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1194 gpio_analog[2] a_289220_348609# a_290737_350685# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1195 a_290737_348985# a_289220_347809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1196 a_5816_240836# a_42877_684772# a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1197 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1198 a_287394_346209# gpio_analog[4] a_287588_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1199 vdda2 a_287812_343783# a_284589_352318# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1200 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1201 a_288222_349659# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1202 gpio_analog[0] gpio_analog[0] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1203 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1204 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1205 a_282219_347336# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1206 gpio_analog[1] gpio_analog[1] vdda1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1207 io_analog[10] a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1208 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1209 a_5816_240836# a_5816_240836# io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1210 vdda1 gpio_analog[1] gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1211 a_42877_684772# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X1212 a_5816_240836# a_287139_344765# a_287144_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1213 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1214 a_540916_680434# a_540916_680434# a_540371_681998# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1215 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1216 a_12801_269626# a_286876_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1217 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1218 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1219 a_288390_344609# a_287350_342628# a_288584_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1220 gpio_analog[2] a_284459_343946# a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1221 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1222 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1223 a_288447_352413# a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1224 a_282219_343936# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1225 a_536916_284434# a_536916_284434# a_290737_348985# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1226 a_287588_346209# a_287812_343783# a_282219_345636# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1227 vdda2 a_287350_342628# a_284589_352318# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1228 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1229 a_24084_271906# a_20532_271136# a_29040_272091# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1230 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1231 gpio_analog[16] a_288222_347259# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1232 gpio_analog[9] a_284459_349046# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1233 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1234 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1235 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1236 io_analog[1] io_analog[1] vccd1 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1237 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1238 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1239 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1240 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1241 a_289220_349409# a_288222_349659# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1242 gpio_analog[9] a_284459_349046# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1243 a_5816_240836# a_20532_271136# a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1244 a_287588_344609# gpio_analog[4] a_287394_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1245 vdda2 a_289220_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1246 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1247 a_290737_350685# gpio_analog[1] a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1248 a_287364_345383# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1249 a_288584_344609# gpio_analog[3] a_288222_344859# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1250 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1251 io_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1252 vdda2 a_287812_343783# a_284689_340388# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1254 a_288222_344059# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1255 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1256 gpio_analog[2] a_289220_349409# a_288447_352413# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1257 a_289220_346209# a_288222_346459# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1258 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1259 a_24084_271906# a_20532_271136# a_29040_272091# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1260 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1261 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1262 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1263 a_540459_681940# io_analog[0] a_540271_687858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1264 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1265 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1266 vdda2 gpio_analog[5] a_287364_345383# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1267 a_5816_240836# a_20532_271136# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1268 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1269 a_5816_240836# a_287139_344765# a_288140_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1270 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1271 vdda2 gpio_analog[4] a_284689_340388# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1272 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1273 a_5816_240836# a_20532_271136# a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1274 a_282219_349036# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 a_5816_240836# gpio_analog[5] a_287364_345383# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1276 a_5816_240836# a_289220_345409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1277 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1278 a_288222_349659# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1279 a_5816_240836# a_284689_340388# a_286876_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1280 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1281 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1282 gpio_analog[2] a_289220_347809# a_290737_348985# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1283 a_289220_343809# a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1284 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1285 a_287812_343783# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 a_288222_346459# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1287 a_288584_348609# gpio_analog[4] a_288390_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1288 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1289 a_40125_693523# a_37693_693523# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X1290 gpio_analog[2] a_284589_352318# gpio_analog[7] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1291 a_5816_240836# a_20532_271136# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1292 vdda2 a_287364_345383# a_284589_352318# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1293 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1294 a_5816_240836# a_42877_684772# a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1295 a_43834_677960# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1296 gpio_analog[2] a_286876_343809# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1297 a_5816_240836# a_288222_344859# a_289220_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1298 a_288390_346209# gpio_analog[5] a_288140_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1299 vccd2 a_43834_677960# a_43834_677960# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1300 a_11871_268125# a_284459_343946# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1301 a_5816_240836# a_5816_240836# gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1302 vdda2 gpio_analog[3] a_288222_348059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1303 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1304 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1305 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1306 vdda1 gpio_analog[0] gpio_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1307 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1308 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1309 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1310 a_5816_240836# a_284589_352318# a_286829_352328# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1311 a_536916_284434# a_536916_284434# a_290737_348985# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1312 vccd1 io_analog[0] io_analog[0] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1313 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1314 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1315 a_287144_346209# a_287364_345383# a_287394_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1316 vdda2 gpio_analog[6] a_287139_344765# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1317 a_5816_240836# a_5816_240836# gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1318 vdda2 gpio_analog[4] a_287350_342628# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1319 gpio_analog[2] a_284459_349046# gpio_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1320 a_540371_681998# a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1321 gpio_analog[12] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1322 gpio_analog[2] a_289220_343809# vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1323 a_5816_240836# a_20532_271136# a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1324 a_288222_344059# a_287364_345383# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 vdda2 gpio_analog[4] a_288222_348059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1326 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1327 a_5816_240836# a_5816_240836# io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1328 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1329 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1330 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1331 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1332 a_290737_348985# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1333 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1334 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1335 vdda2 gpio_analog[6] a_288222_344859# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1336 gpio_analog[8] a_282219_350736# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1337 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1338 a_20532_271136# a_24084_271906# a_24084_271906# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X1339 vdda2 a_282219_347336# a_284459_347346# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1340 gpio_analog[2] a_282219_345636# gpio_analog[11] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1341 a_288447_352413# a_289220_349409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1342 a_288140_344609# a_287364_345383# a_288390_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1343 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1344 gpio_analog[2] a_284459_349046# gpio_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1345 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1346 a_5816_240836# a_5816_240836# gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1347 a_287350_342628# gpio_analog[4] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1348 vdda2 gpio_analog[5] a_284689_340388# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1349 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1350 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1351 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1352 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1353 a_287350_342628# gpio_analog[4] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1354 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1355 a_288447_352413# a_289220_349409# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1356 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1357 gpio_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1358 a_20532_271136# a_284459_342246# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1359 vdda2 gpio_analog[13] gpio_analog[13] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1360 gpio_analog[2] a_289220_345409# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1361 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1362 vdda2 a_288222_348059# a_289220_347809# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1363 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1364 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1365 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1366 a_288222_344859# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1367 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1368 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1369 a_290737_348985# a_289220_347809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1370 io_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1371 gpio_analog[13] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1372 a_284459_342246# a_282219_342236# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1373 vdda2 gpio_analog[6] a_282219_350736# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1374 a_42819_684860# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1375 a_5816_240836# a_541059_678436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1376 a_536459_285940# gpio_analog[0] a_536271_291858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1377 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1378 a_20532_271136# a_284459_342246# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1379 a_12801_269626# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1380 gpio_analog[7] a_284589_352318# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1381 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1382 gpio_analog[2] a_284459_347346# gpio_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1383 a_12801_269626# a_286876_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1384 gpio_analog[2] a_288222_346459# gpio_analog[15] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1385 a_290737_348985# a_289220_347809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1386 a_287394_347809# a_287350_342628# a_287588_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1387 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1388 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1389 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1390 a_288140_347009# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1391 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1392 a_287144_345409# gpio_analog[6] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1393 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1394 vccd1 a_540916_680434# a_540371_681998# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1395 io_analog[9] io_analog[9] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1396 a_12801_269626# a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1397 a_282219_350736# a_287812_343783# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1398 a_290737_348985# a_289220_347809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1399 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1400 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1401 vdda2 a_287364_345383# a_288222_348059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1402 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1403 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1404 a_12801_269626# a_286876_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1405 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1406 a_40125_693523# io_analog[8] a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1407 a_12801_269626# a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X1408 a_29040_272091# a_20532_271136# a_24084_271906# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1409 a_43026_690893# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1410 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1411 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1412 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1413 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1414 a_287588_347809# a_287812_343783# a_282219_349036# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1415 a_40125_693523# a_43026_690893# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1416 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1417 io_analog[10] a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1418 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1419 a_12801_269626# a_286876_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1420 io_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1421 a_288222_347259# gpio_analog[3] a_288584_347009# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1422 a_282219_347336# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1423 a_282219_343936# a_287812_343783# a_287588_345409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1424 a_537154_685355# io_analog[1] a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1425 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1426 gpio_analog[2] a_282219_350736# gpio_analog[8] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1427 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1428 a_20532_271136# a_282219_342236# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1429 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1430 vdda2 a_289220_343809# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1431 a_284459_349046# a_282219_349036# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1432 gpio_analog[2] a_282219_347336# gpio_analog[10] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1433 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1434 a_287812_343783# gpio_analog[3] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1435 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1436 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1437 a_287394_343809# gpio_analog[5] a_287144_343809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1438 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1439 a_290737_350685# gpio_analog[1] a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1440 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1441 a_288447_352413# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1442 gpio_analog[2] a_289220_349409# a_288447_352413# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1443 vdda2 a_287812_343783# a_282219_343936# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1444 a_5816_240836# a_541059_678436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1445 a_288222_345659# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1446 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1447 a_5816_240836# a_5816_240836# gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1448 a_536459_285940# gpio_analog[0] a_536271_291858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1449 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1450 a_5816_240836# a_41723_677112# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1451 a_290737_348985# a_288222_348059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1452 gpio_analog[2] a_288222_349659# a_288447_352413# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1453 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1454 a_540371_681998# a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1455 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1456 a_289220_347809# a_288222_348059# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1457 a_5816_240836# a_5816_240836# io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1458 gpio_analog[12] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1459 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1460 a_5816_240836# a_5816_240836# io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1461 vdda2 gpio_analog[3] a_287812_343783# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 vdda2 gpio_analog[4] a_282219_343936# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1463 a_284589_352318# a_287139_344765# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 gpio_analog[2] a_284459_342246# a_20532_271136# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1465 a_5816_240836# gpio_analog[3] a_287812_343783# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1466 gpio_analog[12] gpio_analog[12] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1467 a_12801_269626# a_284689_340388# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1468 gpio_analog[2] a_288222_348859# a_290737_350685# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1469 gpio_analog[2] a_282219_343936# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1470 a_287394_349409# a_287364_345383# a_287144_349409# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1471 gpio_analog[15] a_288222_346459# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1472 gpio_analog[10] a_284459_347346# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1473 vdda2 gpio_analog[6] a_287139_344765# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1474 a_5816_240836# a_5816_240836# gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1475 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1476 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1477 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1478 a_42819_684860# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1479 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1480 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1481 a_289220_345409# a_288222_345659# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1482 a_43834_677960# a_43834_677960# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1483 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1484 gpio_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1485 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1486 gpio_analog[10] a_284459_347346# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1487 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1488 gpio_analog[2] a_289220_347809# a_290737_348985# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1489 vdda2 gpio_analog[12] gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1490 io_analog[9] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1491 gpio_analog[2] a_289220_344609# gpio_analog[14] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1492 a_5816_240836# a_287139_344765# a_287144_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1493 a_42877_684772# a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.24e+06u l=1e+06u
X1494 vdda2 a_288222_344059# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1495 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1496 a_288390_347809# a_287364_345383# a_288140_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1497 a_288390_346209# a_287350_342628# a_288584_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1498 a_287350_342628# gpio_analog[4] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1499 vdda2 gpio_analog[3] a_288222_349659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1500 a_282219_347336# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1501 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1502 a_11871_268125# gpio_analog[12] a_17579_272227# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1503 gpio_analog[2] a_286876_343809# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1504 gpio_analog[12] gpio_analog[12] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1505 a_5816_240836# gpio_analog[6] a_288140_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1506 gpio_analog[9] a_282219_349036# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1507 vdda1 a_536916_284434# a_290737_348985# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1508 a_540916_680434# a_540371_681998# a_541059_678436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1509 gpio_analog[2] a_282219_342236# a_20532_271136# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1510 a_287144_347809# gpio_analog[5] a_287394_347809# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1511 a_284689_340388# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1512 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1513 a_287588_346209# gpio_analog[4] a_287394_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1514 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1515 a_288222_345659# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1516 gpio_analog[10] a_282219_347336# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1517 vdda2 gpio_analog[4] a_288222_349659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 a_288584_346209# gpio_analog[3] a_288222_346459# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1519 a_5816_240836# gpio_analog[4] a_287350_342628# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1520 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1521 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1522 a_5816_240836# a_288222_345659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1523 gpio_analog[16] a_289220_347009# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1524 vdda2 gpio_analog[12] gpio_analog[12] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1525 vccd1 a_540916_680434# a_540916_680434# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1526 vdda2 a_282219_350736# a_284459_350746# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 gpio_analog[1] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1528 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1529 a_540916_680434# a_540371_681998# a_541059_678436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1530 a_288584_344609# a_287350_342628# a_288390_344609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1531 gpio_analog[2] a_288222_344059# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1532 vdda2 a_287364_345383# a_282219_343936# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1533 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1534 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1535 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1536 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1537 vccd2 a_40125_693523# io_analog[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1538 vdda2 gpio_analog[3] a_288222_344059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1539 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1540 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1541 a_537154_685355# io_analog[1] a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1542 vccd1 a_540271_687858# a_537154_685355# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1543 gpio_analog[12] gpio_analog[12] vdda2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1544 a_20532_271136# a_284459_342246# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1545 io_analog[2] a_540371_681998# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1546 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1547 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1548 a_5816_240836# a_5816_240836# io_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1549 a_290737_350685# a_288222_348859# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1550 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1551 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1552 gpio_analog[2] a_288222_348059# a_290737_348985# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1553 vdda2 a_288222_349659# a_289220_349409# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1554 a_5816_240836# a_537059_282436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=6.9e+07u
X1555 a_5816_240836# a_282219_343936# a_284459_343946# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1556 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1557 a_5816_240836# a_41723_677112# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X1558 gpio_analog[2] a_288222_344859# gpio_analog[14] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1559 vccd2 a_43026_690893# a_43026_690893# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1560 a_540459_681940# io_analog[0] a_540271_687858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1561 vdda1 a_536271_291858# a_290737_350685# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1562 a_17579_272227# a_20532_271136# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1563 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1564 io_analog[8] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1565 a_5816_240836# a_290737_348985# a_536459_285940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1566 a_5816_240836# a_42877_684772# a_42819_684860# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1567 vccd2 a_43026_690893# a_40125_693523# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1568 vdda2 a_287350_342628# a_288222_344059# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 a_5816_240836# a_5816_240836# gpio_analog[1] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1570 gpio_analog[2] a_284459_347346# gpio_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1571 a_288222_348059# gpio_analog[6] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1572 gpio_analog[2] a_284689_340388# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1573 a_536459_285940# gpio_analog[0] a_536271_291858# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1574 a_5816_240836# a_5816_240836# io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1575 a_5816_240836# a_42877_684772# io_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1576 a_530722_289355# a_290737_350685# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=1e+07u
X1577 a_5816_240836# a_288222_346459# a_289220_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1578 a_5816_240836# a_540371_681998# a_540459_681940# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1579 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1580 vdda2 a_14374_271026# a_11871_268125# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1581 vdda2 a_11871_268125# a_12801_269626# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1582 a_287364_345383# gpio_analog[5] vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1583 a_288140_348609# a_287139_344765# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1584 io_analog[10] a_40125_693523# vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1585 a_11871_268125# a_282219_343936# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1586 gpio_analog[2] a_284459_347346# gpio_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1587 a_287364_345383# gpio_analog[5] a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1588 a_5816_240836# a_42877_684772# io_analog[10] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1589 a_11871_268125# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1590 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1591 gpio_analog[2] a_282219_349036# gpio_analog[9] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1592 gpio_analog[11] a_282219_345636# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1593 vdda2 gpio_analog[5] a_288222_349659# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1594 a_12801_269626# a_11871_268125# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1595 vdda1 a_290737_350685# a_288447_352413# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1596 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1597 vdda2 a_288222_344059# a_289220_343809# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1598 io_analog[10] a_42877_684772# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1599 a_5816_240836# a_537059_282436# a_5816_240836# sky130_fd_pr__res_xhigh_po_5p73 w=5.73e+06u l=6.9e+07u
X1600 a_288447_352413# a_288222_349659# gpio_analog[2] vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1601 gpio_analog[14] a_289220_344609# gpio_analog[2] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1602 vccd1 a_540271_687858# a_540271_687858# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1603 vdda2 gpio_analog[5] a_287364_345383# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 vccd2 io_analog[9] io_analog[9] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1605 io_analog[9] a_5816_240836# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1606 vdda2 gpio_analog[6] a_288222_346459# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1607 gpio_analog[2] a_288222_345659# a_5816_240836# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1608 vdda2 a_287139_344765# a_282219_342236# vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 a_290737_348985# a_290737_348985# a_5816_240836# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X1610 gpio_analog[2] a_289220_347009# gpio_analog[16] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1611 a_288222_348859# gpio_analog[3] a_288584_348609# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1612 a_282219_350736# a_287350_342628# vdda2 vdda2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1613 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1614 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1615 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1616 vccd2 io_analog[8] io_analog[8] a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1617 a_5816_240836# a_20532_271136# a_12801_269626# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1618 a_17579_272227# gpio_analog[12] a_11871_268125# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1619 a_288140_346209# gpio_analog[5] a_288390_346209# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1620 io_analog[9] io_analog[9] vccd2 a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X1621 vccd1 a_537154_685355# io_analog[2] vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1622 a_536916_284434# a_290737_348985# a_537059_282436# a_5816_240836# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1623 vccd2 a_43834_677960# a_42877_684772# vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

