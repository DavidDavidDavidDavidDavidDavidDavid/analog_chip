* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_UXPKRJ a_n621_n5174# a_114_n5088# a_n29_n5000# a_n474_n5088#
+ a_n323_n5000# a_461_n5000# a_167_n5000# a_69_n5000# a_16_5022# a_310_n5088# a_n519_n5000#
+ a_n82_n5088# a_n225_n5000# a_363_n5000# a_408_5022# a_212_5022# a_n376_5022# a_n421_n5000#
+ a_n278_n5088# a_n127_n5000# a_265_n5000# a_n180_5022#
X0 a_n421_n5000# a_n474_n5088# a_n519_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X1 a_n225_n5000# a_n278_n5088# a_n323_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X2 a_69_n5000# a_16_5022# a_n29_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X3 a_167_n5000# a_114_n5088# a_69_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=0p ps=0u w=5e+07u l=200000u
X4 a_363_n5000# a_310_n5088# a_265_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X5 a_n29_n5000# a_n82_n5088# a_n127_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=200000u
X6 a_n323_n5000# a_n376_5022# a_n421_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X7 a_n127_n5000# a_n180_5022# a_n225_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X8 a_265_n5000# a_212_5022# a_167_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X9 a_461_n5000# a_408_5022# a_363_n5000# a_n621_n5174# sky130_fd_pr__nfet_01v8 ad=1.45e+13p pd=1.0058e+08u as=0p ps=0u w=5e+07u l=200000u
.ends

.subckt diode_connected_nmos m1_60_4610# m1_120_80# VSUBS
Xsky130_fd_pr__nfet_01v8_UXPKRJ_0 VSUBS m1_120_80# m1_120_80# m1_120_80# m1_60_4610#
+ m1_60_4610# m1_120_80# m1_60_4610# m1_120_80# m1_120_80# m1_60_4610# m1_120_80#
+ m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_120_80# m1_60_4610#
+ m1_60_4610# m1_120_80# sky130_fd_pr__nfet_01v8_UXPKRJ
.ends

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VPWR Y VNB VPB
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=2.05e+12p pd=1.41e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_BDZ9JN a_15_n500# a_n177_n500# a_n561_n500# a_879_n500#
+ a_111_n500# a_n129_n597# a_n513_n597# a_n609_531# a_63_n597# a_n273_n500# a_n801_531#
+ a_687_n500# a_n321_n597# a_159_531# a_639_n597# a_n941_n500# a_783_n500# a_399_n500#
+ a_n81_n500# a_n849_n500# a_351_531# a_n33_531# a_495_n500# a_n897_n597# a_831_n597#
+ a_447_n597# a_n225_531# a_591_n500# a_n657_n500# a_207_n500# a_543_531# a_n753_n500#
+ a_n369_n500# a_303_n500# a_255_n597# a_n705_n597# a_n417_531# w_n1079_n719# a_n465_n500#
+ a_735_531#
X0 a_15_n500# a_n33_531# a_n81_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X1 a_n369_n500# a_n417_531# a_n465_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X2 a_n657_n500# a_n705_n597# a_n753_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X3 a_879_n500# a_831_n597# a_783_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.55e+12p pd=1.062e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X4 a_303_n500# a_255_n597# a_207_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X5 a_n273_n500# a_n321_n597# a_n369_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X6 a_591_n500# a_543_531# a_495_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X7 a_n849_n500# a_n897_n597# a_n941_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.55e+12p ps=1.062e+07u w=5e+06u l=150000u
X8 a_207_n500# a_159_531# a_111_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X9 a_n177_n500# a_n225_531# a_n273_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X10 a_495_n500# a_447_n597# a_399_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X11 a_n561_n500# a_n609_531# a_n657_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X12 a_111_n500# a_63_n597# a_15_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X13 a_783_n500# a_735_531# a_687_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X14 a_399_n500# a_351_531# a_303_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X15 a_n465_n500# a_n513_n597# a_n561_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X16 a_687_n500# a_639_n597# a_591_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X17 a_n753_n500# a_n801_531# a_n849_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X18 a_n81_n500# a_n129_n597# a_n177_n500# w_n1079_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_KBNS5F a_15_n500# a_n177_n500# a_111_n500# a_n273_n500#
+ a_159_n588# a_63_522# a_255_522# a_399_n500# a_n81_n500# a_351_n588# a_n417_n588#
+ a_n129_522# a_n225_n588# a_n321_522# a_n563_n674# a_207_n500# a_n461_n500# a_n369_n500#
+ a_303_n500# a_n33_n588#
X0 a_n81_n500# a_n129_522# a_n177_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X1 a_15_n500# a_n33_n588# a_n81_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X2 a_n369_n500# a_n417_n588# a_n461_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.55e+12p ps=1.062e+07u w=5e+06u l=150000u
X3 a_n273_n500# a_n321_522# a_n369_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X4 a_303_n500# a_255_522# a_207_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X5 a_n177_n500# a_n225_n588# a_n273_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6 a_207_n500# a_159_n588# a_111_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X7 a_111_n500# a_63_522# a_15_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8 a_399_n500# a_351_n588# a_303_n500# a_n563_n674# sky130_fd_pr__nfet_01v8 ad=1.55e+12p pd=1.062e+07u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sized_switch m1_970_n860# m1_1100_n50# m1_1190_n720# m1_3210_n860# w_2760_n990#
+ VSUBS
XXM1 m1_1100_n50# m1_1100_n50# m1_1100_n50# m1_1190_n720# m1_1190_n720# m1_970_n860#
+ m1_970_n860# m1_970_n860# m1_970_n860# m1_1190_n720# m1_970_n860# m1_1190_n720#
+ m1_970_n860# m1_970_n860# m1_970_n860# m1_1100_n50# m1_1100_n50# m1_1100_n50# m1_1190_n720#
+ m1_1190_n720# m1_970_n860# m1_970_n860# m1_1190_n720# m1_970_n860# m1_970_n860#
+ m1_970_n860# m1_970_n860# m1_1100_n50# m1_1190_n720# m1_1100_n50# m1_970_n860# m1_1100_n50#
+ m1_1100_n50# m1_1190_n720# m1_970_n860# m1_970_n860# m1_970_n860# w_2760_n990# m1_1190_n720#
+ m1_970_n860# sky130_fd_pr__pfet_01v8_BDZ9JN
Xsky130_fd_pr__nfet_01v8_KBNS5F_0 m1_1190_n720# m1_1190_n720# m1_1100_n50# m1_1100_n50#
+ m1_3210_n860# m1_3210_n860# m1_3210_n860# m1_1190_n720# m1_1100_n50# m1_3210_n860#
+ m1_3210_n860# m1_3210_n860# m1_3210_n860# m1_3210_n860# VSUBS m1_1190_n720# m1_1100_n50#
+ m1_1190_n720# m1_1100_n50# m1_3210_n860# sky130_fd_pr__nfet_01v8_KBNS5F
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt analog_mux OUT SIG0 SIG1 SIG2 SIG3 SIG4 SIG5 SIG6 SIG7 SIG8 SIG9 SIG10 SIG11
+ SIG12 SIG13 SIG14 SIG15 SEL0 SEL1 SEL2 SEL3 GND VDD
Xx1 x8/A x9/B x9/C x9/D GND VDD x1/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx2 x8/A x9/B x9/C SEL0 GND VDD x2/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx3 x8/A x9/B SEL1 x9/D GND VDD x3/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx4 x8/A x9/B SEL1 SEL0 GND VDD x4/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx5 x8/A SEL2 x9/C x9/D GND VDD x5/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx6 x8/A SEL2 x9/C SEL0 GND VDD x6/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_1 x2/Y OUT SIG1 sky130_fd_sc_hd__inv_2_2/Y VDD GND sized_switch
Xx7 x8/A SEL2 SEL1 x9/D GND VDD x7/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_0 x7/Y OUT SIG6 sky130_fd_sc_hd__inv_2_15/Y VDD GND sized_switch
Xsized_switch_2 x3/Y OUT SIG2 sky130_fd_sc_hd__inv_2_3/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_11 x13/Y GND VDD sky130_fd_sc_hd__inv_2_11/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_10 x12/Y GND VDD sky130_fd_sc_hd__inv_2_10/Y GND VDD sky130_fd_sc_hd__inv_2
Xx8 x8/A SEL2 SEL1 SEL0 GND VDD x8/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsky130_fd_sc_hd__inv_2_12 x14/Y GND VDD sky130_fd_sc_hd__inv_2_12/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_3 x4/Y OUT SIG3 sky130_fd_sc_hd__inv_2_0/Y VDD GND sized_switch
Xx9 SEL3 x9/B x9/C x9/D GND VDD x9/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsky130_fd_sc_hd__inv_2_13 x15/Y GND VDD sky130_fd_sc_hd__inv_2_13/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_4 x5/Y OUT SIG4 sky130_fd_sc_hd__inv_2_5/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_14 x16/Y GND VDD sky130_fd_sc_hd__inv_2_14/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_5 x6/Y OUT SIG5 sky130_fd_sc_hd__inv_2_6/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_0 x4/Y GND VDD sky130_fd_sc_hd__inv_2_0/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_6 x11/Y OUT SIG10 sky130_fd_sc_hd__inv_2_9/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_15 x7/Y GND VDD sky130_fd_sc_hd__inv_2_15/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 x8/Y GND VDD sky130_fd_sc_hd__inv_2_1/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_7 x10/Y OUT SIG9 sky130_fd_sc_hd__inv_2_8/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_2 x2/Y GND VDD sky130_fd_sc_hd__inv_2_2/Y GND VDD sky130_fd_sc_hd__inv_2
Xsized_switch_8 x12/Y OUT SIG11 sky130_fd_sc_hd__inv_2_10/Y VDD GND sized_switch
Xsized_switch_9 x13/Y OUT SIG12 sky130_fd_sc_hd__inv_2_11/Y VDD GND sized_switch
Xsky130_fd_sc_hd__inv_2_3 x3/Y GND VDD sky130_fd_sc_hd__inv_2_3/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_4 x1/Y GND VDD sky130_fd_sc_hd__inv_2_4/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_5 x5/Y GND VDD sky130_fd_sc_hd__inv_2_5/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_6 x6/Y GND VDD sky130_fd_sc_hd__inv_2_6/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_7 x9/Y GND VDD sky130_fd_sc_hd__inv_2_7/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_8 x10/Y GND VDD sky130_fd_sc_hd__inv_2_8/Y GND VDD sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_9 x11/Y GND VDD sky130_fd_sc_hd__inv_2_9/Y GND VDD sky130_fd_sc_hd__inv_2
Xx20 SEL0 GND VDD x9/D GND VDD sky130_fd_sc_hd__inv_8
Xx10 SEL3 x9/B x9/C SEL0 GND VDD x10/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_10 x14/Y OUT SIG13 sky130_fd_sc_hd__inv_2_12/Y VDD GND sized_switch
Xx11 SEL3 x9/B SEL1 x9/D GND VDD x11/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_11 x15/Y OUT SIG14 sky130_fd_sc_hd__inv_2_13/Y VDD GND sized_switch
Xx12 SEL3 x9/B SEL1 SEL0 GND VDD x12/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx13 SEL3 SEL2 x9/C x9/D GND VDD x13/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_12 x8/Y OUT SIG7 sky130_fd_sc_hd__inv_2_1/Y VDD GND sized_switch
Xx15 SEL3 SEL2 SEL1 x9/D GND VDD x15/Y GND VDD sky130_fd_sc_hd__nand4_2
Xx14 SEL3 SEL2 x9/C SEL0 GND VDD x14/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_13 x9/Y OUT SIG8 sky130_fd_sc_hd__inv_2_7/Y VDD GND sized_switch
Xsized_switch_14 x1/Y OUT SIG0 sky130_fd_sc_hd__inv_2_4/Y VDD GND sized_switch
Xx16 SEL3 SEL2 SEL1 SEL0 GND VDD x16/Y GND VDD sky130_fd_sc_hd__nand4_2
Xsized_switch_15 x16/Y OUT SIG15 sky130_fd_sc_hd__inv_2_14/Y VDD GND sized_switch
Xx17 SEL3 GND VDD x8/A GND VDD sky130_fd_sc_hd__inv_8
Xx18 SEL2 GND VDD x9/B GND VDD sky130_fd_sc_hd__inv_8
Xx19 SEL1 GND VDD x9/C GND VDD sky130_fd_sc_hd__inv_8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_95KK7Z c1_n1650_n1600# m3_n1750_n1700#
X0 c1_n1650_n1600# m3_n1750_n1700# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_49C6SK a_n1314_n597# a_524_n500# a_n50_n597# a_n682_n597#
+ a_1156_n500# a_1214_n597# a_n1472_n597# a_682_n500# a_50_n500# a_740_n597# a_1372_n597#
+ a_n840_n597# a_1314_n500# a_n1630_n597# a_840_n500# a_n108_n500# a_1472_n500# a_1530_n597#
+ a_n266_n500# a_n898_n500# a_n1056_n500# a_1630_n500# a_n1688_n500# a_n424_n500#
+ a_108_n597# a_n1214_n500# a_n208_n597# a_n582_n500# a_266_n597# w_n1826_n719# a_208_n500#
+ a_n1372_n500# a_898_n597# a_n366_n597# a_n740_n500# a_424_n597# a_n998_n597# a_n1156_n597#
+ a_366_n500# a_n1530_n500# a_998_n500# a_1056_n597# a_n524_n597# a_582_n597#
X0 a_524_n500# a_424_n597# a_366_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_1630_n500# a_1530_n597# a_1472_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_n1056_n500# a_n1156_n597# a_n1214_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_1156_n500# a_1056_n597# a_998_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_n108_n500# a_n208_n597# a_n266_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_208_n500# a_108_n597# a_50_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1214_n500# a_n1314_n597# a_n1372_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1314_n500# a_1214_n597# a_1156_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X8 a_n740_n500# a_n840_n597# a_n898_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_n582_n500# a_n682_n597# a_n740_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X10 a_682_n500# a_582_n597# a_524_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n266_n500# a_n366_n597# a_n424_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_840_n500# a_740_n597# a_682_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n1530_n500# a_n1630_n597# a_n1688_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_366_n500# a_266_n597# a_208_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_n1372_n500# a_n1472_n597# a_n1530_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_1472_n500# a_1372_n597# a_1314_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_n898_n500# a_n998_n597# a_n1056_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_50_n500# a_n50_n597# a_n108_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_n424_n500# a_n524_n597# a_n582_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 a_998_n500# a_898_n597# a_840_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_JT3SH9 a_1261_n500# a_1319_n588# a_n1319_n500# a_1061_n588#
+ a_n287_n500# a_n1061_n500# a_n1519_n588# a_n487_n588# a_745_n500# a_n1261_n588#
+ a_545_n588# a_1777_n500# a_1577_n588# a_229_n500# a_n1577_n500# a_n545_n500# a_29_n588#
+ a_n1777_n588# a_1003_n500# a_n745_n588# a_803_n588# a_n1937_n674# a_n29_n500# a_487_n500#
+ a_n1835_n500# a_n229_n588# a_n1003_n588# a_287_n588# a_1519_n500# a_n803_n500#
X0 a_n1577_n500# a_n1777_n588# a_n1835_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_1519_n500# a_1319_n588# a_1261_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_n1061_n500# a_n1261_n588# a_n1319_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_1003_n500# a_803_n588# a_745_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_487_n500# a_287_n588# a_229_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_745_n500# a_545_n588# a_487_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 a_1777_n500# a_1577_n588# a_1519_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X7 a_1261_n500# a_1061_n588# a_1003_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 a_n29_n500# a_n229_n588# a_n287_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X9 a_229_n500# a_29_n588# a_n29_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X10 a_n1319_n500# a_n1519_n588# a_n1577_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X11 a_n545_n500# a_n745_n588# a_n803_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X12 a_n803_n500# a_n1003_n588# a_n1061_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 a_n287_n500# a_n487_n588# a_n545_n500# a_n1937_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_F7BMVG a_n573_n1432# a_n703_n1562# a_n573_1000#
X0 a_n573_n1432# a_n573_1000# a_n703_n1562# sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_JEXVB9 a_1261_n500# a_1319_n588# a_n1319_n500# a_1061_n588#
+ a_n287_n500# a_n1061_n500# a_n1519_n588# a_n487_n588# a_745_n500# a_n1261_n588#
+ a_545_n588# a_n1679_n674# a_229_n500# a_n1577_n500# a_n545_n500# a_29_n588# a_1003_n500#
+ a_n745_n588# a_803_n588# a_n29_n500# a_487_n500# a_n229_n588# a_n1003_n588# a_287_n588#
+ a_1519_n500# a_n803_n500#
X0 a_1519_n500# a_1319_n588# a_1261_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_n1061_n500# a_n1261_n588# a_n1319_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_1003_n500# a_803_n588# a_745_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_487_n500# a_287_n588# a_229_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_745_n500# a_545_n588# a_487_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 a_1261_n500# a_1061_n588# a_1003_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 a_n29_n500# a_n229_n588# a_n287_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X7 a_229_n500# a_29_n588# a_n29_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 a_n1319_n500# a_n1519_n588# a_n1577_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X9 a_n545_n500# a_n745_n588# a_n803_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X10 a_n803_n500# a_n1003_n588# a_n1061_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X11 a_n287_n500# a_n487_n588# a_n545_n500# a_n1679_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_9F67JW a_2973_n500# a_n345_n500# a_n1609_n500# w_n3327_n719#
+ a_n1135_n500# a_29_n597# a_n977_n500# a_n2557_n500# a_n129_n597# a_n1767_n500# a_187_n597#
+ a_n503_n500# a_n2083_n500# a_129_n500# a_n1293_n500# a_n287_n597# a_n2715_n500#
+ a_n3031_n500# a_819_n597# a_n1077_n597# a_287_n500# a_n661_n500# a_n1925_n500# a_345_n597#
+ a_n2499_n597# a_n2241_n500# a_n919_n597# a_n1451_n500# a_977_n597# a_n445_n597#
+ a_n2873_n500# a_n1709_n597# a_n2025_n597# a_919_n500# a_2399_n597# a_n1235_n597#
+ a_445_n500# a_503_n597# a_n2657_n597# a_1609_n597# a_n1867_n597# a_n603_n597# a_n2183_n597#
+ a_1077_n500# a_1135_n597# a_661_n597# a_n1393_n597# a_2499_n500# a_2557_n597# a_603_n500#
+ a_2083_n597# a_1767_n597# a_n2815_n597# a_1709_n500# a_1293_n597# a_n761_n597# a_n3131_n597#
+ a_2025_n500# a_n2341_n597# a_1235_n500# a_n1551_n597# a_2657_n500# a_761_n500# a_3031_n597#
+ a_2715_n597# a_n2973_n597# a_2183_n500# a_1867_n500# a_2241_n597# a_1925_n597# a_n29_n500#
+ a_1451_n597# a_1393_n500# a_2873_n597# a_n187_n500# a_3131_n500# a_2815_n500# a_2341_n500#
+ a_n3189_n500# a_1551_n500# a_n2399_n500# a_n819_n500#
X0 a_n661_n500# a_n761_n597# a_n819_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_919_n500# a_819_n597# a_761_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_n187_n500# a_n287_n597# a_n345_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_761_n500# a_661_n597# a_603_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_2025_n500# a_1925_n597# a_1867_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_n2241_n500# a_n2341_n597# a_n2399_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_2341_n500# a_2241_n597# a_2183_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_287_n500# a_187_n597# a_129_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n1293_n500# a_n1393_n597# a_n1451_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_1393_n500# a_1293_n597# a_1235_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_n2873_n500# a_n2973_n597# a_n3031_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X11 a_2973_n500# a_2873_n597# a_2815_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_n345_n500# a_n445_n597# a_n503_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X13 a_n2399_n500# a_n2499_n597# a_n2557_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_2499_n500# a_2399_n597# a_2341_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X15 a_129_n500# a_29_n597# a_n29_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X16 a_1709_n500# a_1609_n597# a_1551_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X17 a_n1609_n500# a_n1709_n597# a_n1767_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X18 a_445_n500# a_345_n597# a_287_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X19 a_n1925_n500# a_n2025_n597# a_n2083_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X20 a_n1451_n500# a_n1551_n597# a_n1609_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X21 a_1551_n500# a_1451_n597# a_1393_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X22 a_n977_n500# a_n1077_n597# a_n1135_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X23 a_n503_n500# a_n603_n597# a_n661_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X24 a_1077_n500# a_977_n597# a_919_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X25 a_n2557_n500# a_n2657_n597# a_n2715_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X26 a_2657_n500# a_2557_n597# a_2499_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X27 a_n29_n500# a_n129_n597# a_n187_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X28 a_603_n500# a_503_n597# a_445_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X29 a_n1135_n500# a_n1235_n597# a_n1293_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X30 a_1235_n500# a_1135_n597# a_1077_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X31 a_n2715_n500# a_n2815_n597# a_n2873_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X32 a_2815_n500# a_2715_n597# a_2657_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X33 a_n3031_n500# a_n3131_n597# a_n3189_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X34 a_3131_n500# a_3031_n597# a_2973_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X35 a_n1767_n500# a_n1867_n597# a_n1925_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X36 a_1867_n500# a_1767_n597# a_1709_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X37 a_n2083_n500# a_n2183_n597# a_n2241_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X38 a_2183_n500# a_2083_n597# a_2025_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X39 a_n819_n500# a_n919_n597# a_n977_n500# w_n3327_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_EJ3ASN a_524_n500# a_108_n588# a_50_n500# a_n208_n588#
+ a_266_n588# a_n366_n588# a_n108_n500# a_424_n588# a_n524_n588# a_n266_n500# a_n50_n588#
+ a_n424_n500# a_n684_n674# a_n582_n500# a_208_n500# a_366_n500#
X0 a_366_n500# a_266_n588# a_208_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n500# a_n50_n588# a_n108_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_n424_n500# a_n524_n588# a_n582_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_524_n500# a_424_n588# a_366_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X4 a_n108_n500# a_n208_n588# a_n266_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_208_n500# a_108_n588# a_50_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X6 a_n266_n500# a_n366_n588# a_n424_n500# a_n684_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_GNAJ57 a_n1314_n597# a_524_n500# a_n50_n597# a_n682_n597#
+ a_1156_n500# a_1214_n597# a_n1472_n597# a_682_n500# a_50_n500# a_740_n597# a_1372_n597#
+ a_n840_n597# a_1314_n500# a_n1630_n597# a_840_n500# a_n108_n500# a_1472_n500# a_1530_n597#
+ a_n266_n500# a_n898_n500# a_n1056_n500# a_1630_n500# a_n1688_n500# a_n424_n500#
+ a_108_n597# a_n1214_n500# a_n208_n597# a_n582_n500# a_266_n597# w_n1826_n719# a_208_n500#
+ a_n1372_n500# a_898_n597# a_n366_n597# a_n740_n500# a_424_n597# a_n998_n597# a_n1156_n597#
+ a_366_n500# a_n1530_n500# a_998_n500# a_1056_n597# a_n524_n597# a_582_n597#
X0 a_524_n500# a_424_n597# a_366_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_1630_n500# a_1530_n597# a_1472_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_n1056_n500# a_n1156_n597# a_n1214_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_1156_n500# a_1056_n597# a_998_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_n108_n500# a_n208_n597# a_n266_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_208_n500# a_108_n597# a_50_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1214_n500# a_n1314_n597# a_n1372_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1314_n500# a_1214_n597# a_1156_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X8 a_n740_n500# a_n840_n597# a_n898_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_n582_n500# a_n682_n597# a_n740_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X10 a_682_n500# a_582_n597# a_524_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n266_n500# a_n366_n597# a_n424_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_840_n500# a_740_n597# a_682_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n1530_n500# a_n1630_n597# a_n1688_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_366_n500# a_266_n597# a_208_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_n1372_n500# a_n1472_n597# a_n1530_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_1472_n500# a_1372_n597# a_1314_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_n898_n500# a_n998_n597# a_n1056_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_50_n500# a_n50_n597# a_n108_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_n424_n500# a_n524_n597# a_n582_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 a_998_n500# a_898_n597# a_840_n500# w_n1826_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt OTA_fingers_031123_NON_FLAT m1_n1130_9530# m1_1130_3110# li_900_7430# m1_n500_70#
+ m1_1130_4630# VSUBS
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_3 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_2 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__pfet_01v8_49C6SK_0 m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730#
+ li_900_7430# m1_90_7730# m1_90_7730# m1_n2620_8810# m1_n2620_8810# m1_90_7730# m1_90_7730#
+ m1_90_7730# m1_n2620_8810# m1_90_7730# li_900_7430# li_900_7430# li_900_7430# m1_90_7730#
+ m1_n2620_8810# m1_n2620_8810# li_900_7430# m1_n2620_8810# li_900_7430# li_900_7430#
+ m1_90_7730# m1_n2620_8810# m1_90_7730# m1_n2620_8810# m1_90_7730# li_900_7430# li_900_7430#
+ li_900_7430# m1_90_7730# m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730# m1_90_7730#
+ m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_90_7730# m1_90_7730# m1_90_7730#
+ sky130_fd_pr__pfet_01v8_49C6SK
Xsky130_fd_pr__nfet_01v8_JT3SH9_0 m1_60_860# m1_n500_70# m1_60_860# m1_n500_70# m1_60_860#
+ VSUBS m1_n500_70# m1_n500_70# m1_60_860# m1_n500_70# m1_n500_70# m1_60_860# m1_n500_70#
+ m1_60_860# VSUBS VSUBS m1_n500_70# m1_n500_70# VSUBS m1_n500_70# m1_n500_70# VSUBS
+ VSUBS VSUBS m1_60_860# m1_n500_70# m1_n500_70# m1_n500_70# VSUBS m1_60_860# sky130_fd_pr__nfet_01v8_JT3SH9
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0 m1_n5940_10010# VSUBS m1_n2620_8810# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1 m1_n5940_10010# VSUBS m1_n2620_8810# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2 m1_n2620_8810# VSUBS m1_n5940_10010# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3 m1_n2620_8810# VSUBS m1_n5940_10010# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__nfet_01v8_JEXVB9_0 VSUBS m1_n500_70# VSUBS m1_n500_70# VSUBS m1_n1130_9530#
+ m1_n500_70# m1_n500_70# VSUBS m1_n500_70# m1_n500_70# VSUBS VSUBS m1_n1130_9530#
+ m1_n1130_9530# m1_n500_70# m1_n1130_9530# m1_n500_70# m1_n500_70# m1_n1130_9530#
+ m1_n1130_9530# m1_n500_70# m1_n500_70# m1_n500_70# m1_n1130_9530# VSUBS sky130_fd_pr__nfet_01v8_JEXVB9
Xsky130_fd_pr__pfet_01v8_9F67JW_0 m1_n1130_9530# li_900_7430# li_900_7430# li_900_7430#
+ m1_n1130_9530# m1_n2620_8810# li_900_7430# li_900_7430# m1_n2620_8810# m1_n1130_9530#
+ m1_n2620_8810# m1_n1130_9530# m1_n1130_9530# m1_n1130_9530# li_900_7430# m1_n2620_8810#
+ m1_n1130_9530# m1_n1130_9530# m1_n2620_8810# m1_n2620_8810# li_900_7430# li_900_7430#
+ li_900_7430# m1_n2620_8810# m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_n1130_9530#
+ m1_n2620_8810# m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_n2620_8810# li_900_7430#
+ m1_n2620_8810# m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# m1_n2620_8810# m1_n2620_8810#
+ m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# m1_n2620_8810#
+ m1_n2620_8810# li_900_7430# m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_n2620_8810#
+ m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# m1_n2620_8810# m1_n2620_8810# m1_n1130_9530#
+ m1_n2620_8810# li_900_7430# m1_n2620_8810# m1_n1130_9530# m1_n1130_9530# m1_n2620_8810#
+ m1_n2620_8810# m1_n2620_8810# li_900_7430# li_900_7430# m1_n2620_8810# m1_n2620_8810#
+ li_900_7430# m1_n2620_8810# m1_n1130_9530# m1_n2620_8810# m1_n1130_9530# li_900_7430#
+ li_900_7430# m1_n1130_9530# li_900_7430# li_900_7430# m1_n1130_9530# m1_n1130_9530#
+ sky130_fd_pr__pfet_01v8_9F67JW
Xsky130_fd_pr__nfet_01v8_EJ3ASN_0 m1_60_860# m1_1130_4630# m1_n2620_8810# m1_1130_4630#
+ m1_1130_4630# m1_1130_4630# m1_60_860# m1_1130_4630# m1_1130_4630# m1_n2620_8810#
+ m1_1130_4630# m1_60_860# VSUBS m1_n2620_8810# m1_60_860# m1_n2620_8810# sky130_fd_pr__nfet_01v8_EJ3ASN
Xsky130_fd_pr__nfet_01v8_EJ3ASN_1 m1_90_7730# m1_1130_3110# m1_60_860# m1_1130_3110#
+ m1_1130_3110# m1_1130_3110# m1_90_7730# m1_1130_3110# m1_1130_3110# m1_60_860# m1_1130_3110#
+ m1_90_7730# VSUBS m1_60_860# m1_90_7730# m1_60_860# sky130_fd_pr__nfet_01v8_EJ3ASN
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_0 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__pfet_01v8_GNAJ57_0 m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730#
+ li_900_7430# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730#
+ m1_90_7730# m1_90_7730# m1_90_7730# li_900_7430# li_900_7430# li_900_7430# m1_90_7730#
+ m1_90_7730# m1_90_7730# li_900_7430# m1_90_7730# li_900_7430# li_900_7430# m1_90_7730#
+ m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# li_900_7430# li_900_7430# li_900_7430#
+ m1_90_7730# m1_90_7730# li_900_7430# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730#
+ m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# m1_90_7730# sky130_fd_pr__pfet_01v8_GNAJ57
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_1 m1_n1130_9530# m1_n5940_10010# sky130_fd_pr__cap_mim_m3_1_95KK7Z
.ends

.subckt constant_gm_local_030423 a_n3719_36# w_n4170_1941# a_n3633_196#
X0 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X1 a_n3688_2136# a_n3688_2136# a_n3633_196# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.348e+07u w=2.5e+06u l=500000u
X2 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=1.74e+13p pd=1.2696e+08u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X3 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X5 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.232e+07u w=1.25e+06u l=1e+06u
X6 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X7 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X9 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X10 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X11 a_n3688_2136# a_n3688_2136# a_n3633_196# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X12 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X14 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X17 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X20 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X21 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X22 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X23 a_n3633_196# a_n3633_196# a_n3719_36# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X24 a_n3688_2136# a_n3633_196# a_n3545_138# a_n3719_36# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X25 w_n4170_1941# a_n3688_2136# a_n3688_2136# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X26 w_n4170_1941# a_n3688_2136# a_n3633_196# w_n4170_1941# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X27 a_n3719_36# a_n3545_138# a_n3719_36# sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_SDAUVS a_n50_n2451# a_n108_n2354# a_n108_118# a_n108_1354#
+ a_n50_1257# a_n50_21# a_n50_4965# a_50_3826# a_50_118# a_50_n3590# a_n50_n1215#
+ a_50_n6062# a_n50_n4923# a_n108_n1118# a_n108_3826# w_n246_n6281# a_n108_n4826#
+ a_n50_n3687# a_n50_3729# a_n50_n6159# a_50_2590# a_50_n2354# a_50_5062# a_n108_2590#
+ a_n108_n3590# a_n50_2493# a_n108_5062# a_n108_n6062# a_50_1354# a_50_n1118# a_50_n4826#
X0 a_50_n6062# a_n50_n6159# a_n108_n6062# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_2590# a_n50_2493# a_n108_2590# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_118# a_n50_21# a_n108_118# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_5062# a_n50_4965# a_n108_5062# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_n4826# a_n50_n4923# a_n108_n4826# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_n2354# a_n50_n2451# a_n108_n2354# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_3826# a_n50_3729# a_n108_3826# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_50_1354# a_n50_1257# a_n108_1354# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_50_n1118# a_n50_n1215# a_n108_n1118# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_50_n3590# a_n50_n3687# a_n108_n3590# w_n246_n6281# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_K6FQWW a_n108_1936# a_n108_n2936# a_n108_718# a_50_n500#
+ a_n50_n3024# a_50_3154# a_n210_n4328# a_50_718# a_n108_n500# a_n50_630# a_n108_n1718#
+ a_n108_3154# a_n108_n4154# a_n50_n588# a_50_n2936# a_n50_1848# a_n50_n1806# a_n50_n4242#
+ a_50_1936# a_50_n1718# a_50_n4154# a_n50_3066#
X0 a_50_n2936# a_n50_n3024# a_n108_n2936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n500# a_n50_n588# a_n108_n500# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_n4154# a_n50_n4242# a_n108_n4154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_1936# a_n50_1848# a_n108_1936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_3154# a_n50_3066# a_n108_3154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_718# a_n50_630# a_n108_718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_n1718# a_n50_n1806# a_n108_n1718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_KG6QWW a_n100_3066# a_n158_1936# a_100_n1718# a_100_n4154#
+ a_100_n500# a_n100_n3024# a_n158_718# a_100_3154# a_n158_n2936# a_n158_n500# a_n158_3154#
+ a_n260_n4328# a_n100_n588# a_n158_n1718# a_n100_1848# a_n158_n4154# a_100_718# a_n100_630#
+ a_100_n2936# a_n100_n4242# a_n100_n1806# a_100_1936#
X0 a_100_718# a_n100_630# a_n158_718# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_100_1936# a_n100_1848# a_n158_1936# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_100_n1718# a_n100_n1806# a_n158_n1718# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_100_3154# a_n100_3066# a_n158_3154# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_100_n2936# a_n100_n3024# a_n158_n2936# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X6 a_100_n4154# a_n100_n4242# a_n158_n4154# a_n260_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_T9YF2H a_n50_n597# w_n246_n4427# a_n108_n2972# a_50_n500#
+ a_n108_736# a_n108_1972# a_n50_1875# a_50_3208# a_n108_n500# a_50_736# a_n50_n1833#
+ a_n50_n4305# a_n108_n1736# a_n108_n4208# a_n50_n3069# a_n108_3208# a_n50_639# a_50_n2972#
+ a_n50_3111# a_50_1972# a_50_n1736# a_50_n4208#
X0 a_50_736# a_n50_639# a_n108_736# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n2972# a_n50_n3069# a_n108_n2972# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_1972# a_n50_1875# a_n108_1972# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_n1736# a_n50_n1833# a_n108_n1736# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_n4208# a_n50_n4305# a_n108_n4208# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_3208# a_n50_3111# a_n108_3208# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_n500# a_n50_n597# a_n108_n500# w_n246_n4427# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_GG6QWW a_100_n3545# a_n100_n2415# a_100_2545# a_n100_n1197#
+ a_n158_n1109# a_n100_1239# a_n100_21# a_n260_n3719# a_100_109# a_n158_2545# a_100_n2327#
+ a_100_1327# a_n158_n3545# a_n158_1327# a_100_n1109# a_n100_n3633# a_n158_109# a_n158_n2327#
+ a_n100_2457#
X0 a_100_1327# a_n100_1239# a_n158_1327# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_100_2545# a_n100_2457# a_n158_2545# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_100_n1109# a_n100_n1197# a_n158_n1109# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_100_n2327# a_n100_n2415# a_n158_n2327# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_100_n3545# a_n100_n3633# a_n158_n3545# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_100_109# a_n100_21# a_n158_109# a_n260_n3719# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_R8BLL7 a_n108_1936# a_n108_n2936# a_n108_718# a_50_n500#
+ a_n50_n3024# a_50_3154# a_n210_n4328# a_50_718# a_n108_n500# a_n50_630# a_n108_n1718#
+ a_n108_3154# a_n108_n4154# a_n50_n588# a_50_n2936# a_n50_1848# a_n50_n1806# a_n50_n4242#
+ a_50_1936# a_50_n1718# a_50_n4154# a_n50_3066#
X0 a_50_n2936# a_n50_n3024# a_n108_n2936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_50_n500# a_n50_n588# a_n108_n500# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X2 a_50_n4154# a_n50_n4242# a_n108_n4154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_50_1936# a_n50_1848# a_n108_1936# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_50_3154# a_n50_3066# a_n108_3154# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_50_718# a_n50_630# a_n108_718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_50_n1718# a_n50_n1806# a_n108_n1718# a_n210_n4328# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt ota_3_11_23_nonflat m1_n6050_3760# m1_n4180_2590# m1_n4190_3090# m1_n4200_780#
+ w_n6280_3640# VSUBS
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_3 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_2 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__pfet_01v8_SDAUVS_0 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__pfet_01v8_SDAUVS_1 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__pfet_01v8_SDAUVS_2 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__pfet_01v8_SDAUVS_3 m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760# m1_n6050_3760#
+ m1_n7530_3520# m1_n6050_3760# m1_n7530_3520# w_n6280_3640# w_n6280_3640# w_n6280_3640#
+ w_n6280_3640# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n6050_3760# m1_n6050_3760#
+ m1_n6050_3760# w_n6280_3640# w_n6280_3640# m1_n7530_3520# w_n6280_3640# w_n6280_3640#
+ m1_n6050_3760# m1_n6050_3760# m1_n6050_3760# sky130_fd_pr__pfet_01v8_SDAUVS
Xsky130_fd_pr__nfet_01v8_K6FQWW_0 m1_n4120_60# m1_n4120_60# m1_n4120_60# m1_n4300_8710#
+ m1_n4180_2590# m1_n4300_8710# VSUBS m1_n4300_8710# m1_n4120_60# m1_n4180_2590# m1_n4120_60#
+ m1_n4120_60# m1_n4120_60# m1_n4180_2590# m1_n4300_8710# m1_n4180_2590# m1_n4180_2590#
+ m1_n4180_2590# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4180_2590# sky130_fd_pr__nfet_01v8_K6FQWW
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0 m1_n7530_3520# VSUBS m1_n9960_3530# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1 m1_n7530_3520# VSUBS m1_n9960_3530# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__nfet_01v8_KG6QWW_0 m1_n4200_780# VSUBS m1_n4120_60# m1_n4120_60# m1_n4120_60#
+ m1_n4200_780# VSUBS m1_n4120_60# VSUBS VSUBS VSUBS VSUBS m1_n4200_780# VSUBS m1_n4200_780#
+ VSUBS m1_n4120_60# m1_n4200_780# m1_n4120_60# m1_n4200_780# m1_n4200_780# m1_n4120_60#
+ sky130_fd_pr__nfet_01v8_KG6QWW
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2 m1_n9960_3530# VSUBS m1_n7530_3520# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__nfet_01v8_KG6QWW_1 m1_n4200_780# VSUBS m1_n4120_60# m1_n4120_60# m1_n4120_60#
+ m1_n4200_780# VSUBS m1_n4120_60# VSUBS VSUBS VSUBS VSUBS m1_n4200_780# VSUBS m1_n4200_780#
+ VSUBS m1_n4120_60# m1_n4200_780# m1_n4120_60# m1_n4200_780# m1_n4200_780# m1_n4120_60#
+ sky130_fd_pr__nfet_01v8_KG6QWW
Xsky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3 m1_n9960_3530# VSUBS m1_n7530_3520# sky130_fd_pr__res_xhigh_po_5p73_F7BMVG
Xsky130_fd_pr__pfet_01v8_T9YF2H_0 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n7530_3520#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n7530_3520# w_n6280_3640# m1_n7530_3520#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n7530_3520# m1_n4300_8710# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_1 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n4300_8710# w_n6280_3640# m1_n4300_8710#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_2 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n7530_3520#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n7530_3520# w_n6280_3640# m1_n7530_3520#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n7530_3520# m1_n4300_8710# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_3 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n4300_8710# w_n6280_3640# m1_n4300_8710#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_5 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n7530_3520#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n7530_3520# w_n6280_3640# m1_n7530_3520#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n7530_3520# m1_n4300_8710# m1_n7530_3520# m1_n7530_3520# m1_n7530_3520#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__pfet_01v8_T9YF2H_4 m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710#
+ w_n6280_3640# w_n6280_3640# m1_n4300_8710# m1_n4300_8710# w_n6280_3640# m1_n4300_8710#
+ m1_n4300_8710# m1_n4300_8710# w_n6280_3640# w_n6280_3640# m1_n4300_8710# w_n6280_3640#
+ m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710# m1_n4300_8710#
+ sky130_fd_pr__pfet_01v8_T9YF2H
Xsky130_fd_pr__nfet_01v8_GG6QWW_0 VSUBS m1_n4200_780# VSUBS m1_n4200_780# m1_n6050_3760#
+ m1_n4200_780# m1_n4200_780# VSUBS VSUBS m1_n6050_3760# VSUBS VSUBS m1_n6050_3760#
+ m1_n6050_3760# VSUBS m1_n4200_780# m1_n6050_3760# m1_n6050_3760# m1_n4200_780# sky130_fd_pr__nfet_01v8_GG6QWW
Xsky130_fd_pr__nfet_01v8_R8BLL7_0 m1_n7530_3520# m1_n7530_3520# m1_n7530_3520# m1_n4120_60#
+ m1_n4190_3090# m1_n4120_60# VSUBS m1_n4120_60# m1_n7530_3520# m1_n4190_3090# m1_n7530_3520#
+ m1_n7530_3520# m1_n7530_3520# m1_n4190_3090# m1_n4120_60# m1_n4190_3090# m1_n4190_3090#
+ m1_n4190_3090# m1_n4120_60# m1_n4120_60# m1_n4120_60# m1_n4190_3090# sky130_fd_pr__nfet_01v8_R8BLL7
Xsky130_fd_pr__nfet_01v8_GG6QWW_1 VSUBS m1_n4200_780# VSUBS m1_n4200_780# m1_n6050_3760#
+ m1_n4200_780# m1_n4200_780# VSUBS VSUBS m1_n6050_3760# VSUBS VSUBS m1_n6050_3760#
+ m1_n6050_3760# VSUBS m1_n4200_780# m1_n6050_3760# m1_n6050_3760# m1_n4200_780# sky130_fd_pr__nfet_01v8_GG6QWW
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_0 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
Xsky130_fd_pr__cap_mim_m3_1_95KK7Z_1 m1_n6050_3760# m1_n9960_3530# sky130_fd_pr__cap_mim_m3_1_95KK7Z
.ends

.subckt OTA_MULT_GM ota_3_11_23_nonflat_0/w_n6280_3640# ota_3_11_23_nonflat_0/m1_n4180_2590#
+ ota_3_11_23_nonflat_0/m1_n4190_3090# constant_gm_local_030423_0/w_n4170_1941# ota_3_11_23_nonflat_0/m1_n6050_3760#
+ VSUBS
Xconstant_gm_local_030423_0 VSUBS constant_gm_local_030423_0/w_n4170_1941# m1_n200_1910#
+ constant_gm_local_030423
Xota_3_11_23_nonflat_0 ota_3_11_23_nonflat_0/m1_n6050_3760# ota_3_11_23_nonflat_0/m1_n4180_2590#
+ ota_3_11_23_nonflat_0/m1_n4190_3090# m1_n200_1910# ota_3_11_23_nonflat_0/w_n6280_3640#
+ VSUBS ota_3_11_23_nonflat
.ends

.subckt sky130_fd_pr__nfet_01v8_A5635U a_229_n125# a_n647_n299# a_n545_n125# a_n487_n213#
+ a_487_n125# a_n29_n125# a_29_n213# a_n287_n125# a_n229_n213# a_287_n213#
X0 a_n287_n125# a_n487_n213# a_n545_n125# a_n647_n299# sky130_fd_pr__nfet_01v8 ad=3.625e+11p pd=3.08e+06u as=3.625e+11p ps=3.08e+06u w=1.25e+06u l=1e+06u
X1 a_487_n125# a_287_n213# a_229_n125# a_n647_n299# sky130_fd_pr__nfet_01v8 ad=3.625e+11p pd=3.08e+06u as=3.625e+11p ps=3.08e+06u w=1.25e+06u l=1e+06u
X2 a_n29_n125# a_n229_n213# a_n287_n125# a_n647_n299# sky130_fd_pr__nfet_01v8 ad=3.625e+11p pd=3.08e+06u as=0p ps=0u w=1.25e+06u l=1e+06u
X3 a_229_n125# a_29_n213# a_n29_n125# a_n647_n299# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_H7FLKU a_29_n338# a_n29_n250# a_n129_n338# a_n187_n250#
+ a_n289_n424# a_129_n250#
X0 a_129_n250# a_29_n338# a_n29_n250# a_n289_n424# sky130_fd_pr__nfet_01v8 ad=7.25e+11p pd=5.58e+06u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=500000u
X1 a_n29_n250# a_n129_n338# a_n187_n250# a_n289_n424# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=500000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_B5N4SD a_n573_6900# a_n573_n7332# VSUBS
X0 a_n573_n7332# a_n573_6900# VSUBS sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_LK874N a_29_n597# a_n287_n500# a_n745_n597# a_745_n500#
+ a_n229_n597# a_287_n597# a_229_n500# a_n545_n500# w_n941_n719# a_n487_n597# a_n29_n500#
+ a_545_n597# a_487_n500# a_n803_n500#
X0 a_n29_n500# a_n229_n597# a_n287_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_229_n500# a_29_n597# a_n29_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X2 a_n545_n500# a_n745_n597# a_n803_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_n287_n500# a_n487_n597# a_n545_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 a_745_n500# a_545_n597# a_487_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_487_n500# a_287_n597# a_229_n500# w_n941_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_GLZPWL a_n287_n500# a_n487_n588# a_745_n500# a_545_n588#
+ a_229_n500# a_n545_n500# a_29_n588# a_n745_n588# a_n29_n500# a_487_n500# a_n229_n588#
+ a_n905_n674# a_287_n588# a_n803_n500#
X0 a_487_n500# a_287_n588# a_229_n500# a_n905_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_745_n500# a_545_n588# a_487_n500# a_n905_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X2 a_n29_n500# a_n229_n588# a_n287_n500# a_n905_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_229_n500# a_29_n588# a_n29_n500# a_n905_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 a_n545_n500# a_n745_n588# a_n803_n500# a_n905_n674# sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_n287_n500# a_n487_n588# a_n545_n500# a_n905_n674# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt constant_gm_fingers Vout VDD VSS
Xsky130_fd_pr__nfet_01v8_A5635U_0 Vout VSS VSS Vout VSS VSS Vout Vout Vout Vout sky130_fd_pr__nfet_01v8_A5635U
Xsky130_fd_pr__nfet_01v8_H7FLKU_0 m1_n210_n170# Vout m1_n210_n170# m1_n210_n170# VSS
+ m1_n210_n170# sky130_fd_pr__nfet_01v8_H7FLKU
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_0 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_1 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_2 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__res_xhigh_po_5p73_B5N4SD_3 m1_n1220_n5790# VSS VSS sky130_fd_pr__res_xhigh_po_5p73_B5N4SD
Xsky130_fd_pr__pfet_01v8_LK874N_0 m1_n210_n170# VDD m1_n210_n170# VDD m1_n210_n170#
+ m1_n210_n170# VDD Vout VDD m1_n210_n170# Vout m1_n210_n170# Vout VDD sky130_fd_pr__pfet_01v8_LK874N
Xsky130_fd_pr__pfet_01v8_LK874N_1 m1_n210_n170# VDD m1_n210_n170# VDD m1_n210_n170#
+ m1_n210_n170# VDD m1_n210_n170# VDD m1_n210_n170# m1_n210_n170# m1_n210_n170# m1_n210_n170#
+ VDD sky130_fd_pr__pfet_01v8_LK874N
Xsky130_fd_pr__nfet_01v8_GLZPWL_0 m1_n210_n170# Vout m1_n210_n170# Vout m1_n210_n170#
+ m1_n1220_n5790# Vout Vout m1_n1220_n5790# m1_n1220_n5790# Vout VSS Vout m1_n210_n170#
+ sky130_fd_pr__nfet_01v8_GLZPWL
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i vdda2 vdda1
Xdiode_connected_nmos_6 vccd1 io_analog[0] analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_7 io_analog[0] analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
Xanalog_mux_0 gpio_analog[2] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_analog[10]
+ gpio_analog[11] analog_mux_0/SIG5 analog_mux_0/SIG6 analog_mux_0/SIG7 vdda2 gpio_analog[14]
+ analog_mux_0/GND gpio_analog[15] gpio_analog[16] analog_mux_0/SIG13 analog_mux_0/SIG14
+ analog_mux_0/SIG15 analog_mux_0/SEL0 analog_mux_0/SEL1 analog_mux_0/SEL2 analog_mux_0/SEL3
+ analog_mux_0/GND vdda2 analog_mux
XOTA_fingers_031123_NON_FLAT_0 io_analog[10] io_analog[9] vccd2 constant_gm_fingers_0/Vout
+ io_analog[8] analog_mux_0/GND OTA_fingers_031123_NON_FLAT
Xdiode_connected_nmos_0 vccd2 io_analog[9] analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_1 io_analog[9] analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_2 io_analog[8] analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
Xdiode_connected_nmos_4 io_analog[1] analog_mux_0/GND analog_mux_0/GND diode_connected_nmos
XOTA_MULT_GM_0 vccd1 io_analog[0] io_analog[1] vccd1 io_analog[2] analog_mux_0/GND
+ OTA_MULT_GM
Xdiode_connected_nmos_3 vccd2 io_analog[8] analog_mux_0/GND diode_connected_nmos
Xconstant_gm_fingers_0 constant_gm_fingers_0/Vout vccd2 analog_mux_0/GND constant_gm_fingers
Xdiode_connected_nmos_5 vccd1 io_analog[1] analog_mux_0/GND diode_connected_nmos
R0 vssd2 analog_mux_0/GND sky130_fd_pr__res_generic_m3 w=7.55e+07u l=1e+07u
X0 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=3.235e+13p pd=2.2294e+08u as=1.3679e+14p ps=1.00302e+09u w=5e+06u l=500000u
X1 a_24084_271906# a_24084_271906# analog_mux_0/SIG6 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=7.25e+12p pd=5.348e+07u as=9.6e+12p ps=6.5e+07u w=2.5e+06u l=500000u
X2 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=7.17999e+14p pd=5.06914e+09u as=4.06e+13p ps=2.9624e+08u w=5e+06u l=1e+06u
X3 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=1.363e+14p pd=9.9452e+08u as=3.045e+13p ps=2.2218e+08u w=5e+06u l=500000u
X4 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.54e+13p ps=3.1816e+08u w=5e+06u l=500000u
X5 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X6 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.595e+13p ps=1.1638e+08u w=5e+06u l=500000u
X7 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=2.555e+13p pd=1.8022e+08u as=0p ps=0u w=5e+06u l=1e+06u
X8 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X9 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.83e+13p ps=1.2732e+08u w=5e+06u l=1e+06u
X10 analog_mux_0/GND analog_mux_0/SIG6 a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+13p ps=1.6928e+08u w=5e+06u l=1e+06u
X11 gpio_analog[13] gpio_analog[13] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=3.18606e+14p ps=2.87548e+09u w=5e+07u l=200000u
X12 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+13p ps=5.2976e+08u w=5e+06u l=500000u
X13 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X14 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X16 vdda2 gpio_analog[13] gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X17 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X21 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X22 gpio_analog[13] gpio_analog[13] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X23 analog_mux_0/GND analog_mux_0/GND gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X24 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X25 vdda1 a_536916_284434# analog_mux_0/SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.51e+13p ps=1.7004e+08u w=5e+06u l=1e+06u
X26 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.685e+13p ps=3.2874e+08u w=5e+06u l=500000u
X27 gpio_analog[12] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
R1 vssa2 analog_mux_0/GND sky130_fd_pr__res_generic_m3 w=7.45e+07u l=2.6e+06u
X28 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X29 analog_mux_0/SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X30 analog_mux_0/GND analog_mux_0/GND gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X31 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X32 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X33 analog_mux_0/GND analog_mux_0/GND gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X34 analog_mux_0/SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X35 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X36 a_17579_272227# gpio_analog[12] analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.395e+13p ps=9.558e+07u w=5e+06u l=500000u
X37 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X38 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X39 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X40 a_530722_289355# analog_mux_0/SIG14 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X41 gpio_analog[12] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X42 vdda2 a_24084_271906# analog_mux_0/SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.075e+13p ps=1.383e+08u w=5e+06u l=1e+06u
X43 gpio_analog[13] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X44 gpio_analog[12] gpio_analog[12] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X45 analog_mux_0/GND analog_mux_0/GND gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X46 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X47 vdda2 gpio_analog[13] gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X48 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X49 gpio_analog[13] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X50 analog_mux_0/SIG5 gpio_analog[12] a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X51 a_536916_284434# analog_mux_0/SIG13 a_537059_282436# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.015e+13p pd=7.464e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=1e+06u
X52 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X53 vdda1 a_536916_284434# analog_mux_0/SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X54 gpio_analog[13] gpio_analog[13] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X55 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X56 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X57 analog_mux_0/GND analog_mux_0/GND gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X58 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X59 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X60 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.105e+13p pd=7.674e+07u as=0p ps=0u w=1.25e+06u l=1e+06u
X61 vdda1 gpio_analog[1] gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=3.81686e+14p pd=3.65032e+09u as=1.595e+14p ps=1.10638e+09u w=5e+07u l=200000u
X62 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X63 a_17579_272227# gpio_analog[12] analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X64 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X65 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X66 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X67 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X68 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X69 gpio_analog[1] gpio_analog[1] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X70 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X71 vdda2 gpio_analog[12] gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X72 a_17579_272227# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X73 gpio_analog[0] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.595e+14p pd=1.10638e+09u as=0p ps=0u w=5e+07u l=200000u
X74 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X75 gpio_analog[12] gpio_analog[12] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X76 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X77 a_17579_272227# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X78 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X79 analog_mux_0/SIG14 gpio_analog[1] a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=1.83e+13p pd=1.2732e+08u as=0p ps=0u w=5e+06u l=500000u
X80 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X81 a_17579_272227# gpio_analog[12] analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X82 vdda2 gpio_analog[12] gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X83 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X84 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X85 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X86 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X87 a_29040_272091# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.72e+06u l=6.9e+07u
X88 vdda1 gpio_analog[1] gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X89 analog_mux_0/SIG6 a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X90 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X91 gpio_analog[1] gpio_analog[1] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X92 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X93 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X94 a_24084_271906# analog_mux_0/SIG6 a_29040_272091# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=1e+06u
X95 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X96 vdda1 a_536916_284434# analog_mux_0/SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X97 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X98 analog_mux_0/SIG5 gpio_analog[12] a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X99 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X100 a_17579_272227# gpio_analog[13] a_14374_271026# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.232e+07u w=5e+06u l=500000u
X101 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X102 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X103 a_536459_285940# gpio_analog[0] a_536271_291858# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.015e+13p ps=7.406e+07u w=5e+06u l=500000u
X104 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X105 analog_mux_0/GND a_537059_282436# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X106 gpio_analog[13] gpio_analog[13] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X107 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X108 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X109 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X110 analog_mux_0/GND analog_mux_0/GND gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X111 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X112 analog_mux_0/GND analog_mux_0/SIG6 a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X113 vdda2 gpio_analog[13] gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X114 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X115 vdda1 gpio_analog[0] gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X116 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X117 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X118 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X119 gpio_analog[13] gpio_analog[13] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X120 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X121 analog_mux_0/GND analog_mux_0/SIG6 a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X122 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X123 analog_mux_0/SIG14 gpio_analog[1] a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X124 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X125 vdda2 gpio_analog[13] gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X126 a_536459_285940# gpio_analog[0] a_536271_291858# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X127 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X128 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X129 analog_mux_0/GND a_537059_282436# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X130 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X131 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X132 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X133 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X134 a_14374_271026# gpio_analog[13] a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X135 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X136 vdda2 a_24084_271906# analog_mux_0/SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X137 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X138 gpio_analog[13] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X139 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X140 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X141 analog_mux_0/SIG14 gpio_analog[1] a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X142 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X143 analog_mux_0/GND analog_mux_0/GND gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X144 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X145 gpio_analog[1] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X146 analog_mux_0/GND analog_mux_0/GND gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X147 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X148 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X149 analog_mux_0/SIG14 a_530722_289355# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X150 gpio_analog[13] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X151 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X152 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X153 gpio_analog[0] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X154 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X155 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X156 analog_mux_0/GND analog_mux_0/GND gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X157 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X158 a_29040_272091# analog_mux_0/SIG6 a_24084_271906# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X159 analog_mux_0/GND analog_mux_0/GND gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X160 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X161 a_29040_272091# analog_mux_0/SIG6 a_24084_271906# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X162 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X163 gpio_analog[0] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X164 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X165 a_17579_272227# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X166 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X167 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X169 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X170 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X171 analog_mux_0/SIG6 a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X172 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X173 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X174 a_14374_271026# gpio_analog[13] a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X175 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X176 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X177 analog_mux_0/SIG14 gpio_analog[1] a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X178 analog_mux_0/GND analog_mux_0/GND gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X179 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X180 gpio_analog[1] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X181 a_536459_285940# gpio_analog[0] a_536271_291858# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X182 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X183 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X185 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X186 a_17579_272227# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X187 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X188 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X189 analog_mux_0/SIG5 a_11871_265693# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X190 analog_mux_0/GND analog_mux_0/GND gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X191 a_17579_272227# gpio_analog[13] a_14374_271026# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X192 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X193 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X194 a_11871_265693# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
R2 analog_mux_0/GND vssd1 sky130_fd_pr__res_generic_m3 w=7.7e+07u l=5e+06u
X195 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X196 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X197 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X198 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X199 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X200 a_14374_271026# gpio_analog[13] a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X201 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X202 vdda1 a_536916_284434# analog_mux_0/SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X203 analog_mux_0/SIG14 a_530722_289355# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X204 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X205 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X206 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X207 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X208 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X209 vdda1 a_536916_284434# analog_mux_0/SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X210 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X211 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X213 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X214 analog_mux_0/GND analog_mux_0/SIG6 a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X215 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X216 analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X217 a_14374_271026# gpio_analog[13] a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X218 gpio_analog[0] gpio_analog[0] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X219 a_536916_284434# analog_mux_0/SIG13 a_537059_282436# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X220 vdda1 gpio_analog[0] gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X221 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X222 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X223 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X224 a_536916_284434# analog_mux_0/SIG13 a_537059_282436# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X225 gpio_analog[0] gpio_analog[0] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X226 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X227 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X228 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X229 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X230 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X231 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X232 vdda1 gpio_analog[0] gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X233 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X234 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X235 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X236 a_29040_272091# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.72e+06u l=6.9e+07u
X237 analog_mux_0/SIG5 a_11871_265693# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X238 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X239 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X240 gpio_analog[0] gpio_analog[0] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X241 a_11871_265693# analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X242 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X243 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X244 analog_mux_0/SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X245 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X246 a_536916_284434# analog_mux_0/SIG13 a_537059_282436# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X247 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X248 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X249 a_17579_272227# gpio_analog[13] a_14374_271026# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X250 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X251 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X252 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X253 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X254 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X255 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X256 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X257 gpio_analog[1] gpio_analog[1] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X258 analog_mux_0/GND analog_mux_0/GND gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X259 vdda2 a_24084_271906# analog_mux_0/SIG6 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X260 gpio_analog[0] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X261 gpio_analog[12] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X262 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X263 vdda1 gpio_analog[1] gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X264 a_29040_272091# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.72e+06u l=6.9e+07u
X265 analog_mux_0/GND analog_mux_0/GND gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X266 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X267 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X268 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X269 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X270 gpio_analog[0] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X271 analog_mux_0/SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X272 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X273 a_17579_272227# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
R3 analog_mux_0/GND vssa1 sky130_fd_pr__res_generic_m4 w=2.75e+07u l=2.8e+06u
X274 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X275 a_536916_284434# analog_mux_0/SIG13 a_537059_282436# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X276 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG6 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X277 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X278 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X279 vdda2 gpio_analog[12] gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X280 a_29040_272091# analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.72e+06u l=6.9e+07u
X281 gpio_analog[1] gpio_analog[1] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X282 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X283 a_17579_272227# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X284 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X285 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X286 analog_mux_0/SIG6 a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X287 analog_mux_0/SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X288 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X289 vdda1 gpio_analog[1] gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X290 vdda2 a_24084_271906# a_24084_271906# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X291 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X292 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X293 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X294 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X295 gpio_analog[0] gpio_analog[0] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X296 analog_mux_0/SIG14 gpio_analog[1] a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X297 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X298 a_536459_285940# gpio_analog[0] a_536271_291858# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X299 vdda1 gpio_analog[0] gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X300 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X301 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X302 gpio_analog[0] gpio_analog[0] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X303 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X304 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X305 gpio_analog[1] gpio_analog[1] vdda1 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X306 vdda1 gpio_analog[1] gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X307 analog_mux_0/SIG15 a_530722_289355# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X308 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X309 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X310 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X311 a_536916_284434# a_536916_284434# analog_mux_0/SIG13 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X312 a_24084_271906# analog_mux_0/SIG6 a_29040_272091# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X313 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X314 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X315 analog_mux_0/GND analog_mux_0/SIG6 a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X316 analog_mux_0/SIG14 gpio_analog[1] a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X317 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X318 a_24084_271906# analog_mux_0/SIG6 a_29040_272091# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X319 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X320 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X321 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X322 a_24084_271906# a_24084_271906# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X323 analog_mux_0/GND analog_mux_0/SIG6 a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X324 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X325 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X326 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X327 analog_mux_0/GND analog_mux_0/GND gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X328 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X329 vdda1 gpio_analog[0] gpio_analog[0] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X330 a_536916_284434# a_536916_284434# analog_mux_0/SIG13 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X331 analog_mux_0/GND analog_mux_0/GND gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X332 gpio_analog[12] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X333 analog_mux_0/GND analog_mux_0/SIG6 a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X334 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X335 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X336 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X337 analog_mux_0/SIG6 a_24084_271906# a_24084_271906# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X338 analog_mux_0/GND analog_mux_0/GND gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X339 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X340 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X341 gpio_analog[1] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X342 vdda2 gpio_analog[13] gpio_analog[13] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X343 gpio_analog[13] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X344 a_536459_285940# gpio_analog[0] a_536271_291858# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X345 analog_mux_0/SIG7 analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X346 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X347 analog_mux_0/SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X348 vdda2 a_14374_271026# a_14374_271026# vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X349 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X350 a_29040_272091# analog_mux_0/SIG6 a_24084_271906# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X351 analog_mux_0/SIG7 a_11871_265693# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X352 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X353 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X354 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X355 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X356 analog_mux_0/SIG14 gpio_analog[1] a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X357 analog_mux_0/SIG15 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X358 analog_mux_0/GND analog_mux_0/GND gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X359 a_536459_285940# gpio_analog[0] a_536271_291858# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X360 gpio_analog[12] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X361 gpio_analog[12] gpio_analog[12] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X362 analog_mux_0/GND analog_mux_0/GND gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X363 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X364 gpio_analog[1] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X365 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X366 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X367 vdda2 gpio_analog[12] gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X368 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X369 analog_mux_0/SIG5 gpio_analog[12] a_17579_272227# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X370 gpio_analog[12] gpio_analog[12] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X371 vdda1 a_536916_284434# analog_mux_0/SIG13 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X372 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X373 vdda2 gpio_analog[12] gpio_analog[12] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X374 gpio_analog[1] analog_mux_0/GND analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X375 gpio_analog[12] gpio_analog[12] vdda2 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X376 analog_mux_0/GND a_537059_282436# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X377 a_17579_272227# analog_mux_0/SIG6 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X378 vdda1 a_536271_291858# analog_mux_0/SIG14 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X379 analog_mux_0/GND analog_mux_0/SIG13 a_536459_285940# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X380 analog_mux_0/GND analog_mux_0/GND gpio_analog[1] analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=200000u
X381 a_536459_285940# gpio_analog[0] a_536271_291858# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X382 a_530722_289355# analog_mux_0/SIG14 analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=1e+07u
X383 vdda2 a_14374_271026# analog_mux_0/SIG5 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X384 vdda2 analog_mux_0/SIG5 analog_mux_0/SIG7 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X385 a_14374_271026# a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X386 analog_mux_0/SIG5 a_14374_271026# vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X387 analog_mux_0/SIG7 analog_mux_0/SIG5 vdda2 vdda2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X388 vdda1 analog_mux_0/SIG14 analog_mux_0/SIG15 vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X389 analog_mux_0/GND a_537059_282436# analog_mux_0/GND sky130_fd_pr__res_xhigh_po w=5.73e+06u l=6.9e+07u
X390 analog_mux_0/SIG13 analog_mux_0/SIG13 analog_mux_0/GND analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X391 vdda1 a_536271_291858# a_536271_291858# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X392 analog_mux_0/GND analog_mux_0/SIG6 analog_mux_0/SIG7 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X393 vdda1 a_536916_284434# a_536916_284434# vdda1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X394 a_17579_272227# gpio_analog[12] analog_mux_0/SIG5 analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X395 a_536916_284434# analog_mux_0/SIG13 a_537059_282436# analog_mux_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

